`timescale 1 ns/1 ns
module ahb2pvci(
	pvci_addr, pvci_wd, pvci_valid, pvci_rd, pvci_rdata,
        hclk, hresetn, haddr, htrans, hwrite, hsize, hburst,
	hsel, hwdata, hrdata, hresp, hready);
//parameter declaration
//**************************************
// input ports
//**************************************	
 //AHB ports	
	input         hclk; 			 // clock
	input         hresetn;			 // active low reset
	input [31:0]  hwdata;			 // data bus		
	input         hwrite;			 // write/read enable
	input [2:0]   hburst;			 // burst type
	input [2:0]   hsize;			 // data size
	input [1:0]   htrans;			 // type of transfer
	input         hsel;			 // slave select 
	input [31:0]  haddr;
  //PVCI ports
        input [7:0]   pvci_rdata;
//**************************************
// output ports
//**************************************
  //PVCI ports
        output [7:0]  pvci_addr;						
        output [7:0]  pvci_wd;
        output        pvci_valid;
        output        pvci_rd;
   
		
 // AHB ports
	output [31:0] hrdata;			 // data output for wishbone slave
	output [1:0]  hresp;			 // response signal from slave
	output        hready;			 // slave ready
`pragma protect begin_protected
`pragma protect author = "MED"
`pragma protect author_info = "VirtuaLAB"
`pragma protect encrypt_agent = "RTLC VELOCE", encrypt_agent_info = "1.5"
`pragma protect key_keyowner = "Mentor Graphics Corporation"
`pragma protect key_keyname =  "MGC-VERIF-SIM-RSA-1"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype =  "base64")
`pragma protect key_block
HJybrNnYyEzTX3OE2urotFPeJ9qtLkZnIW8S2jJbktQP5UdwIt3jVpvGK+OZDcc4
5OuNBnqasP0/x2BnQbE4VyIJYka3yzh3htJ3Cvtmd42LASlMyapv8tTwqCOtBPdJ
jreYiCQlxQvUFfRFgYnnIvv2AJSS/exLgwIejHD2zAY=
`pragma protect key_keyowner = "Mentor Graphics Corporation"
`pragma protect key_keyname =  "MGC-VELOCE-RSA"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype =  "base64")
`pragma protect key_block
luGr1ugTYMox4DVNdm+h0QEGeTmxLiCwHO3y13ofMV/vVC1+G7/LJ3OQAorV0Vvn
03vIYHm77+pz6xJiomTHQbWumQJwYwS6eESzhKtsZ+e41ozY5JIyP1gSRisSf64P
jSEwKXdGYERMP8q5L7QpB85is58eWsmN0BH/1spxo9E=
`pragma protect data_method =  "aes128-cbc"
`pragma protect encoding = ( enctype =  "base64" )
`pragma protect data_block
xEGECptdpCIMrOEAfEyaIfzzHJUitq/5zLxmRqjfOGgZr4FweiiaiTWUnLMI0nmv
hWYavOPWQEMa6+1cOtb5eh1QBbhsUZH3k5bwbZq2GlCk1mbTlJGVGo4WEmQCBfhu
l+6jqc4f0bOV6Nk5LQyv3bta2OeHDNChoJABuaYBRpCn2STeBA6YhDbPbcXAEKrj
enhPHfTHx8BZn2CcUUnSbTlDo69dgvf/FlZydD/lEnE8oMBA1+r9W8K3gjpGuk1j
gbTVdO9V/2i+lnTptde9thRlz+RJRXKMvuVF/Ny/yymlVRvGOfiS5TaeHBty9K6m
xLN9LlkPUhRaDYDU115rpDccB6mpIYH35t8vWivPqZVs+Hsp6C1TVI92hOGKhBsJ
TzHrDC2dFPWlOAahGEB9aQpozoJSJh+9EdFIW8PG/zpED3vj7JtERWp5wGmuROR9
kI2GtdVV7MXh4VZS57t1xwvFtuI6a4KRjbBWFpQbjzO4neGc+tfZ6A89pMZG9k8h
TQnS2FLatcBaNiss19D3PjYW5NopDv4seksejXoB2CAnFYO7OHs4Jq4KFunb/DFo
7FtptDv6/QsuN3Gtyy4Q9xhRdN2HOpL+e0jAUnX4PUTeY6CKBwiQdnrrB0NPaGff
0chIvu0zPC7M5tOT1Ht3yrN5TbA29nwmj7JuA6eTNWV1DwK7k9hx/lccHU5tywdM
2rXWMOn83EoLGer0k6U6Vncxogw6qUrFUjuKhba0CaoCMlFJzLG7O8Qc7ub9WHv0
CzBFqJksnTJrRfDFStlZSKqfDKvyiBqVczSyo/j2ezSIGFNkrPqQq3cap4ABTyf5
GgqE2oDk8WInPZEemVxkp/L6R9+BdvocyubJTzh53eTR7Z8BOgTuRmgXQYRa2gwr
icog140WqquhZFiwVESLepOGSPentPNjLP5GmCVB+oaEyLuOOmwlYZ+OiAGUDkC5
Oq/iFAVJv95abKd6V4Ukg7mVWbmtl91CtmnUb5pE2eXPuLLvZgFhSWgtd0u+m/9s
gKMHIkMXkWYTQyx1WXLwViGviAA0BOcIVBpSWt+jVvRtaTj0L9MxUU/StWjDKUaD
FiuDdSjzL8x0YWF8T+tmHvXGxIJx1Qw/+PJegdw45leIYT2RqvFHPivB0ZsgJnl4
2eQtPDa/sWxcF08WMw6+P/xywCggl2yjzXnxNxRNNhsROg1xCpgGF3ZluQWUnXWz
T8ayMHL3tOQq3O2OWdca3sDtTxDpUAhFcR+5BLHDeL/ewCpsWaaHPn7G8t0OO5+O
FaC0WCNmK88kHGu1DZkUueQY39MTP4p3nfpbHQRQMoCJp5bqivi23+DlWmo1OkIJ
RUEMCZwIEpX2fp/gc+8EnSrNIFALwOXDs4gzIUh25PqehDfXXiBu1oz3YbuCgQLZ
vUTU6f4IVnaOvGr0xFv5+X2E5jOYH+4h73IU336/Po54XX1KzkNtE6z/soaMW+UB
8w3Q0Jf8oobvP3TywB1/2KzFAaCPlXkIrecMzw0/bh0mZB1y/HnlTMS3Da7K7DX7
MJQMO/ABwfGuj248D8pgw0EDItiBDAXvzkNgCqE51z72VI+P/maKLs+rFvd7vxt6
YVIw129WF6nVs+nVT83P2ufD+h/TqE6yb28CGW/wVLbVRSU1jcUAYsMp4TfxrARn
6Ruxn6vk8kVQTN9px1ddcWtP+h2n5ijeMJIpviMsV3ZWhD8tSPG3f37Vhh6sRdVh
A50Oq7FYSOAqab1RMCabXR+FKj4/Ea1Pjd2MnasM0my3+AOUCM2qB1B12ZKp/pW5
gRbcJC/JhGqPRhNSKbGjTA0sBahASRImE4+0HO9rxp9gC0UtDksC3UPwBVCqXwho
QyKN11Bc+SvLiArsHs/O6kj7WqpWE3R0lCYAZIR/4H+GNOWXLvTc4p6GW2SThqT8
R9FIaF+gVy2vsRpy9Nj6HgF1GsNjfklzRB7UOjMzoTY24E/UtHqVdM7vXqb4DV2C
yYsORveSt/8OYKdslbOewRH+kwC8OZ1QVQfaM5miwVD4H1jT5QUKUUGEgWhNwzdp
EOfFknLynitl/TrBZLpDallnt4lyIdkpa7Bq805Ql40W/kEKfB16Qgp2eHp9LByw
vBaQwzdVydOWEinawWymSqFAmXZLWbmMprrcLFBwDcP61S8N1/xJt8hypFduBZE0
Px6aFaKJo/2ZEbjXKtl6Hd4UwJms3LkIMriLin2fFClrYi47Zm9623TwettRD7fR
W7/yYj7PxL8OqUqT47scola+vGDmSUd6Qdrr+lO98Tg+m+8Kxbm7omdqWuchNPy5
U2FUj4Kw6FUfley85/X0LOVAz4HvGrp609LZnUHjHgBIqTrt83Q6Bw3gjhdCHhqE
C+v3+kYySM5+4BMElIefboHXDL07fsFe9T93g4x4g1Ylm7wsc0bmigkgTvVYYxDI
Xh2boiVN+mLIS7R1xpXt/afdyNYYtc4DZApykKo24IZEoaJDO7oCDZWxIfjoFSrJ
9f7b09lG+Z6lLd3f59i/ZYHQTm97Hni825BomDjY/fLYnxFXJIUrsBrNSeD6fu5m
88jGcpjzLQyBPLTops5NVeDWxl8JTUXXmoiWT9Z2skXU3pdI0yVjnRc13vjSNe9E
SfTQKcVXh6HArDTRl8owxf+6E9X2iTcDG97I7v+4J/d8NOVIQafGJ2L8SN246sae
Rs5mKKF0echE0wMJQSXXo3AmMwCAGfFlNqgUY6vP5w178f1lqMrEy43d9HTib9P9
fjM/Uxm9uqV2QHcy0RDd50Dpe4CNBCv+sEAX2CRZ36lHpnku4wqmW2C4DQXhGJTz
2GUYR3BVIBGiVXHxiHgErcXFytGjJ+5UiM2S4H7rAJRPSQ2rAXwR4TRz4OUDt5Sx
Y+o/N1t2yJ5WnzcuJVrnLC1esjQJ0WbLCwuH4ieMAHNzs2lkI3e1JY9qmyGU76zL
gGMGwKaf5KpP0rzwd+BzZhZ9cVwbWGwo7PVDYOVyAXLFNQ+ujfnc+vbZVFUg91/H
6CTQ5c9jPRd5tqxJCuAbsBqb60gohfeJKvWFvIYx0VEz3N3WvW21SHRfGcBfH2Ql
FdQp/ekumsXyF2fq2abXUIgKQm+16Oup8LxC1q0g9jxbSZ3/85DvN5H5/zIHq8Ae
x4QvxGW89g/CGUd/mfhwKs0WS5fZ8KVTMheligFpWogyzDEgDrDsk8oAi/W1Pmai
8G9d/meC/I7NZsXlWi9x9/6I+0tpUxAHjgpsKmr19igIeknG+lYv5qkOPuvaP3IU
GkNCSEUVzGBvMzMPZKqfqI1NC2YdoRYX5RO/GxcM5MYgfp/JUx4ibXBV8/QaQ+2t
3vX2qTNGF9JLlgCcKsaHJ9UR+tpu6GGEfO9mY4tZu3HhwVp3/fBmU6qvUbDDB69r
VGm1wUwoMhwWQFSeN8/dWUCB2gYh5xyR7VnS1t/Ci1NRjxzm7SoeQUIUM1H5lxWA
jarQicHKJd1iMkNBKXUez+rouCII40y4PrBMcU5ytzxfRtzLTIdU5eOtrB4BNEdD
5g+dKywzS1NBlZOklgTiTMJrmOM0CdMpDUgba3mZTFLd5twh5BteQNVDTnX8cbDx
xrVovRSGL3Wz+3NqHCnkCGAz0KQjl5kHwv9NAZItdQ+yGdI/7Ubt2Sj73b0K/t9o
11q87fPPMf2/C3VWS6oGqAHyuCMBRe/5WKPgJNUW6rwlnZbeXGJs0UdtzILEcjxn
G690w7WO4pLlVBsVp2bE0WeXkbTC0HMJ54R7h7T38eet4Jts/hZYxAsv/VyAU4pm
ulhYLb3sK21n2gAXKncCDBwd3zMA9JdDCP5FIcfdT0HFHnmO6dE0LgNRP7+fqxyj
Hak/qL2S8CidhC4VFpxu6a0479v2cz5G39rEgrjvZ3rgDOBvf+ipfVkrhmsRrAD8
lRikA5UmY0QGZOMyfyyTP/C3W+6kL9DUXor1TDlJl+eYqAe54IYi3xOGMyh56GFD
iop530bB7RVdMWGxICsnmz2rr4c8mEeQBzhrEpu95AyV/Co7BqBoEmteX0Gf8lTe
b8qXYNOyKExCAwW4aizUgQRTOz1L6e4UsQuKLvMuj8HovUXG8NqKwo+T7O5zfExq
uWZ4Nzv4gaXYyGdHmFUVlYA+i7XbkLvXo++/y459HjzT6msn2AFQNnxha9DC247M
CM+LrguHF/kLp9kOCiviQU43oZ3Yk/F8ZIe/FB71RBt8RgOJCfxcUAy8LvxnuH3/
YC8wvAqezTsq+/C49V8Ft2kmMD/VwggNAtURKE+iwyDvGxDi95iVKxIY5Bgf2qOS
opq0XJcyYB0IaRusuJyJGmkvJ2N3nRfkkkqfbW69rdlLjbNYBkLy42RzrzLBtr9i
f0WDFChXxzDO8soxQrcfUFnfmtbAb/9kWjyrrQyUC72H5g2XWF816XK17lVMaxTO
lpany7a0yT2bIyOKkmvwltee/wkq0UCXROAaOAu4KlCriCVaHbMsqHBdGULszeC6
DHbv/4C44mPuey3ZFaVKhabYFMDwSyST0uIImcRyagu72pflwuy98g69D9PWOzKs
gH4qBLCamTEJR8SaUbHNiWor4f3d4CBuNm1/gwWVruObrc81pKXlYa2oie2sOaLj
71zQjVtU+qCv6iDvGPQUBnfyaju7Z2ipUhwzgyTsXK4g+RCv4QkyA/yXobKPRS/B
Oz8Xk/7pKm2x3hJaFybdODc4LwieZqUT7ibq3UkS1kpmXjQXevuVSjOi6NC3Y2XA
vmAUUz1bcabunGW3dOd33J7tMPP87igKfnJls7w97C/MjWk8Xw+rlf38+MnEYKhW
wvb6QWIcp8hwiv4ShmptN0gm4+3aZTOL8tzfXN7+pgdnAd4iWsGeGXTm2mWU3qQs
l+Z1GoBwhCRQtAWOTGHtO9f7tViEbMRglCuv5Q18PUvQuRju3emvO+l22fKyZD1y
I18mAu6n99DOQFUxCWMwBCjAUHOkEPoUdFdoVmA10y6OMRi8qEoLCFM7eTscOjeP
XEjaYiQyFngu8S3RzAL4o7Gfccv+Y8Dv36mYXIUTj2wrTIUNHBk4uPNCYgIsnOSj
1ko97aAQ2OQEAuwdFXIEeMjl4e+JDuHJc6Tkv014dfEK6u/w4DfSYVxJbwS92T4f
MY3TitRI0DmbjlDf84mUmWv2/Km+o/dQHuUYDr+HVq4MP/ggyjw2olSasLhK3cuy
2k//09kBF7t3YNTCYTIFnpbEmGx0XdXnUnE+c69RGV9NfHUUFhYTgGeKZxxlnpGt
h1yFlClmabSndAUUpUF+bGhs+/dDuELWdn7pF+EAFHHS9lEmddFpsAmbPwsFgiu/
bVAX1cyG6xpCEnVhV7gTM1zMcimvfg/ziQbweJwDri3qL/eLnO0X2P7oBv09aig5
yETQFTTuKwzklVbZeqRZZ7iSrxrWS9oVWs5fkF8+zKcqXXf9f1Mv2ThGkaQ8NJx9
U/ZDUP7ZI5XTlI7FXk3kaq0rCdbpeN0fzOfnNtJNNl6tXUJttLamelhTXiEx7JRF
hL94IaUHwNArjnh2XNnTf40kWmnBWOA7JXUb5EWz6kK1krEeP+HC65y5SyPjr3RW
mJf6HU/lBw9z5txp4vTWWoyxtA/pWkRUovVRSd3vDmGTI1Z+2mmNSbgJgvaFiW9u
vjM7+90EJOMt5o+Q1xXTv1KGLEdd2K5CIjvUnZuWVnSFRWhi5rt+WHvl5zcBD11V
wHpBZwJtpya/nfp3YRTrj7LhlQl99DU2TfNfjiq9ddm0Ua2RedM9zBI9QYq0haz0
rLcZzRRld4UNzyengQmush1stUPYGm5LmEPMB4E/zoNUhBylLw9hBaMgEcaX9cno
bcwFxkoFtucKg0eEI16czJ8pl7qdSqVNdTm6uV++Lc7PsoGFYMCKIEd9kVx6FY3q
s0y5iCWW2oJli6noejplvESgl9Wt+SxAGCHFR/UW9VAg7nAvYwy41ynozBJIsT9H
t23AP4i8bhk+OEiGXowD+F+ODAZMWzxBlsHPDNJYMFruppYpo7xZNAf2HbjMRPen
g0YAK6tpzenRJvmr5Sn/BuYnRNJwUmlybsVuR/BjC2im4eggiuRwM7qpoHfoveI6
NxwyGnLxWMvVh42lC9I4I+Zkys3fPu4f9Vv9iHcSRCaEKcWIC+I62uzmLP/IAZ+v
FjIAzNVHMDF39TipkqwMIwlU1fGiRW2ihkMMCx6xr1pLeKcS2suCN6vHOoOCvzM3
Rhtq1GpuVzKPxoYpIYdOaq5sG2XQDpF8sm9rDEroMC11oi4+jo61wx1FWzYYTuyI
8gHYvqS8w5M16loF2N3FZ15O3cQijRASgEfNWmVcWHyDHAIAkYA2CW5N4EtRSCgQ
ecVVEVzbK4vNrQ0T5Inj+/A+e2hNy3azDQd4DtctI+TpOAjSKuLvkiTr/90A2y8p
Nz4gBTEvK7Mbn/SNvkQAvIpg86hTT6JPquWEG/D29mqJUaXBaX3uKwmlHufGnbn9
mEW4DobvAH8GaAUHKDhQ5MIrMbtNTNZGh3K/a1TLaEttKtBWqWYpIgRfdyoJFU3p
rDIIYTO8cWj0s3Kvw3P2fq9X4rVPJdskqNu5LCcMpB7G8HDqoAFFexH3CLDrjp/B
934MYDArm8S2dkSBH8AkDEsi6oLxOjGdWQMBtTEkEBmi1QKRNgcdedzugBRB6YLs
mzg4mP99Y+gE0qC1yOk4n1UfSUFzZVXRHgq7B+TgrqAthTgbMBSStW1/7xtQbRJQ
YTtjr06Ly+x9sAFYOUOSpW301jARY2uKH8qqhK333R91sm0HGlBw/qtwDXVrUPdf
IToFM/mPaBOjqTtAy3mvMkBwMjbuSCEt9i78Ly+RZu4T/JRjbg2NWZAb/x8l+doS
pVTsyHx+n4v+LmPHgo8RU0d04N6T4hmaGkUmufs6miQiWpIyrF6DLoYsNewOvaU3
sD2wy6lC77A1Mq/sS2sMByCcyUFc3tx8OT2N7biABLShhxx9vS+zuVSvOMpsYzDv
IfCK1fIeW95RzVz1QRYZSxZUvse8EffbLgMCNEoM2YYMhk+yDL/Bv1jdyfNAMBJY
lI7ipXTZFN/HUGTVSjSe4kVMC8quVakjhgwszIjdHCa1h1gs3FanpJhjypPyauKT
C4O/p0OoCzMi4vay+IYa1dmXQ0BtNASAf3ZgH7M7WhTN+vTDczTJRjH6cEULbM4m
o9ASNRweeU/b6+CXssGJ2FVDOaLQG5/opckr0aM7qVgdx5P7rTHRJZOloAHR3SF7
Ip416yCmb3QvpgVB7EjvPPEiy32ZPosRjd3JEXRNb7qsKXHam02QRvzbXZJuZqlk
P3I88GUkbwCG6p7bjqnrz6mgSmibYH3u/REU/BEKHg5WCRph2SZL7hLnV7O5V3y5
cxy0k3QfEZ1i0b0xAbl6GttXcDYb07VpO6owzVJaqvKOp2rctyPc+mhZ/RNcfWGI
v0hNgX8r205F3Y8u2Dy+Wymd7+uiAlvulPq+6oBsYgkphCylK3vRWr0hayTeSCQa
9wSj4h6kKMyCs+sE6c0jOb7krCPXQsnO8ONY1T7sM257pUsRadkO09O3tGcDL/U2
ohcJxW33pPTuGS6xLYVCCKbJU/yvolxR7TjXF2B7neTh42on5bE5fd/8apZoRG1q
vqS7hXhePdwSVIyaZ5lPTcmBt4MFzXn8cO+/sPoiyRq7OG9m1/FUypsXVg44Vpm7
LJCqqcDr7Zk8JQ8g0YWB5TYrgN863CBk5mVifBtHtT0E4FLrMPq5fS2cCZyNg7BV
i1eCv/95wN2U21tOweIFMbrP2IpnEbgQkW6gtQXX4Buw3U6y2xCIc9gvgXccKz3d
4vOSYPgfW7hQZ5khSD1hQI/cD6uagFXlRQeUK0ZEWJixM/UKqyM4bk59WUi1/lwF
3qJQS/xz8tDS8VfdMG6imMSqnoggL1ORVxjtboDl55xfKYtVYeJ1vYy0x9WcLeXD
kXnpT1KEAjaJOn+xyhhyQq0k8hgc8qNOm+LT1jh5TStwuRnR4CCFoknO7zIV0QuD
NBLPeKqIjAAFoAxAxBQFzWXPe1Cs/xe9NKGFCS85YRPwfqzevlPdAG9vix18Xdy2
+jBXnaGiYpWSlkvFt+ZbOS/9xljJO6G2XoqDxN/Vyi8cllnvgQvCesYOcYqwlgz/
ZgKXItG+RbwREj96rTFJ6bdbHxFdNCJb1zKuBYXzqdQ3tMWOqRttr9S8tNxbr2D1
18NFcJ+icMolaWySFmXN/sSs109nZxRrS/SemUlFa576BlETD59xf5Caz4gt6hcg
lSjHlPijvK2+2WiJ2s/HDyHJdwZnowXJ/vJK01g6XzwFdNo+UNGStC7jD9kupRPj
rOz4nz0uz3pj695RwA4TVEnUFHGxpN77s6AoNT+Lc8gjs2dusg4YfBLKaXDPh6kx
HfnQ6A/R2VKYraGQos338cy/Kbe1SpC+7Si1sp2lXt7JBhGPbS60XynfYkEhObNK
vHMs9sbp4Ygcq2b7qA2nNXT0U0qoIi4GqahmUHp7eHf3Zga/uQMLhzOMzF8qDXId
W3jQCsr22B61dmS2/3Wpcxg4+MYUeVaAQs2AeHWDYUl/JUnwXZ3RXUI4SuM8XX7e
VXhI6d6zRqfSZfK+INrMJWHJfH7EXOig3qNuKk1i3V6Ca543jQMyl+jHG5bRXYBZ
rDE9PmynN/XpWPKhoSpbC0a3x1orBGPRMl8zfDHl/dvgJAg1fgRazeiu/io2asmL
Tpn/9l0TiX7dpyae70nF3K3JnNjiLpJJXChjNLShK9Co8CEte+56ZxqLhQWpmJ5T
zsrjfU1slnHZ0l4PA6Fm5bmqWsbvlPQZAcMGMAlOJgmjG8757U1an1kFQiAw0oQT
iPnUAqcO+v8Jj+8brPbPzZrO/+Iy8PuUnp3H1bD9uKcg8R8Iv4k2EglPsKipG2xt
Nb6IUy723ZorO/uWdtRcZebl61ldtv4+RnvH1k3XNWSuLs5F1sZ+ro0Pc/drOT7Z
o21HkNgjdjAOv/dkZpBHK1UT8abtg3O2+2PQdsfLYj7sykfqyJC0UqFYibQx3ejf
KU5xoehZ7zXaZPw4dR7hzlpWzXdcurVmxlSJsjsdX2Prou4YD1e8ET6aDjFbtOay
MulUBgtNc66f0kbyIybAToUH3hqQbgArvNh5jjDU+9PgLAL+pFyLzsZ+9MtDCSak
rnmpcogwlgiUx0KCxTn09Nq+DubiuPvDp4o30EcJ5YIrGp5p1rno6aNOWNzaXRRB
tUOVE+o/ZZLbDmelvQ7pqZV1kL8Q0QwiVMuwybKur9814k0QXhrYhJi7yoOc7bEH
0WsfpV8/UZLvp1anyQmm5Yn0NT2TYHhDVAewaeUyQmltLT8rcfqSzO43fUxgtDWU
PIyhLZDhVhc7bqE3FpWxhRun75wfhw/bLQ/zDGFGfdRST+iu+8wN43QpoQHjX9w2
r7jVjZs4nSZWMWoCnvgbuRD0T0EfvL4d5NsgXyS/H3XE0ccnGxRzxjCh6Z/ovybt
R28HyIEdSPaq7XXAHNp7eDcCQ3U5Yb0zwIlMqrndFPLlKWRc0zQcsogSPyqXO+4R
MmyCkps5tl6iJA9IdZDRWtvFYlG7YhWuJ+m4RQXZ8J6g5M0PlZ5a4PBf8Q1PknSE
F2kRiFSUC3Cmt6RyWdGSkcU1JIw98SrrMAn3xG1RLqY5msYwjlocYpU1zvSFKGmj
G0PWvmrBPBMv/KLXJbPnioKClpa/McqzBKPRofehwaWLFrzTp+gJ5tbRNtFP+m9q
UEREdLiEogahwzqKzG2LgwxsXRxZiJIkXoHam5fsorLgNozvjwRVpwYeHBOoEFnT
RFGIexxnc7n65EXccIORPamoixJiqLJhTRRT/Ux6tFmq9bQ2Hud6pOZYqq+qyrLl
pFy44uY1FW3mmtpMijA7pWY4hKLXIcshzD3yIYwehUBK/ZuVPvBkuCoJ6jY+ScVe
/pWrSEoATecMczlohpmiEWuo/P9QwkM0bf3eBAQEFDUkTQkxtoz4aIjSD5hETOSY
5AGX34ty8K2f1BpwlWIWBhRKWv2MqEibu2kwufPS9xX1FzszaLSJ70VGMPJ5Kz4Q
FG1av48ILjYo1bywXcBJNXS1m4FCOeHK1owt8hDqQ4F3pwlVw95z4MDsY/BvDNWc
W4mMLNgQvClclWCZkbj0/SujX9ou01qXbj20HfYUSGVFDY8sZaJR5+lBQVrf6kZ3
3Qekt+DMNc5ryjL5g+fzyOjKq5swZOjFMdelvu9cp39DwiXLzjnW7wXSBVGYPlfp
EjL0XbmCXIi10aDatbxdhu/bC4qrucYa8qDHRSWtOlgds/2f4oGxY3IS1ZP2yQpC
C/S9zA8eqfnD5lHfvHAmtpa9SAMP2vR9nqdB0LXWR3DaheafwA+SeLoVFyGGbFCo
w4cLaRn+/XPc/K3DtUrAVCx6Y1rIexCp3mUtqybDs34GG0trSMyQYLw5kLDxX6rK
JUTcWz3aEIYLyVQcQEJzJYYZ+mBZaJcb//93CKuzEoVqfPiECNqDMx9vutdnl0PL
aZ1UfcguOOX/dbuOQ40snFmqsraeBtLXSxokIlhDhEje0bxa2wYCo/FgkOA9bHcy
VMkPbRAMh7AJrVD1P4KR+3Nlawwp3D09me6hcXNKCJm2J8dQn/etNUkRMRIEamEc
nkjNSGTLvqVopPwN3r0pe9UJCKMvnV6poeB3IEU/tSAonlJCTBLdhd4DCkgepmOk
tlaMMeIEZnCrCEEu+sjBUkW9SbK47Xsp+y1p5qFHPOwRzLygvOkMYDbIMOp3aENt
xFwF7zJUXMGTDUqijg1NATNBWdt84tcImOZT5McvAx0k+xon11N+uFkVmMPqW/vX
CqZBW7jU83XRkrNUxwAXIN9IvyIH+n8enN+2tRwC8CwdIgn6FJ35nwEVv6Zm1Gb2
vShXM94xcR8ZyOTkpzEpZZJpSRWfllgeAvvrJrqTjYRqaqJ0++3D1yOy22CLYnMS
abW4HN5yNdYBsQqn3EpiHlf8EwYg4WcFo7rtIsgcbBoLTq59MnBaUxegqQ2ctKLg
zHgSLMZ3VZAPEFziEpr1ghSA/eiZ0k+ocpntwB+KURUXpbKOJ4QPYOif36Hpwl2s
gjQBHGXyjd3nJkOGbJTufFQ+gKE7tB02zE+ayxPPStk18xuNXdu4PPf82CZdG5TX
5ouxZ2j8kAMmsGdbR7H+9xyhckrWaeh8yXk9JvVFkmESzUUg445Ocq3/CoTmiX+J
GUcRUCEk0KzQ8CLsj1kifEcPQ4g/zK4JA0K9eZcEJSAWo9+URLwil+Kb7kBaju0O
0lFDpVTcZOJKtZ3IZ53s99gVIPUHXo+8ho5irZ3IWRdW1Z4N0F0fa+W6pNbzO5FA
P3z7oLVdvY5vyKKga/MLa4P1k93mjZj3rN1UoPFH/8hmkDCIJ67MOtFuv4QGmOtF
8/X8j93aK9W1tn3aRvCf0pPpVkyDZ2Yt71b+dOiMOWIAMwMzDOOG5SlPnfEE36f3
nOV6AZBN4sY50Yegel4+sI7zpMkluBFU3jMQhrs05dFiBak6N0bpzvooB+NWZZCl
CibBIkp4qZ8UaRahUiskQF5UpHLyXPeETW50uBgbnEz9192MJGaKLhvbWGIBWnVl
cfgnJmw0U2WHtw0rVfSl3soGQjjSav91HWVM5i0NhBDQGcqpGupC8KJC9X1Jt9A3
87iy7ozmFg8qfpVZb9Cdl6D7LWybdh9+dDbAe5PCP7TIaNyck5TdskrYNnDJnR6s
eeOjy/xrXhacp0sGtxz+8YDTgz9cqyD6EJ7/ynuiki4l7WU8XCPuaw2ddoqiXZJL
AHMtYptDQhuRk3ihKLi1fcjKiA9YafczN+zMOtI00t1lDMDOkUmAuEYLtXyZTY4o
/zaFezrtYxhzBW27hm3kuI++JapbWZsK5umXEykskS/kFauO/3y4rokTMWXDtXUi
400nxMmm6U9igVmD+zufIB2fDjP4hHSIwMYdTuBuwOyysV90dxu15GSbhBcKoTly
bFBAvUqs45NY5UUDac+XeF88jOd9FmQggTgWnoej514dPWQBcu+lAJi30b9s0vve
mdAZhBi/ELjSWfq3KOdmapebGFovWwFBkM5x5QZZ48H43gD98655FocU+mdbrLYB
CPOhwO4erEmMOBYGWaXwdVytarAHGP3xoWlsQy7Q3q39+0cobbYt6QGcCaNHpt9n
be5vT3y3T6zhoajq4EpBkstiP+8+sOt9VlduCITd5eEG1BJ0lVOWWIdAoTqZiGwi
83xnSruKz4B4MQp54gASQDRNZR/qwSYJbA7LRTjbrT9Fr+ht8n4xWCEhnM0oO/6m
C/c4OoEaVYpzT5nXse2Tf395cnfRzfQXapBTJOfXCwU2o4VwXnFiEFu7G50JLzgi
6gS4SkmqwWrCwjnj82bxzdwbshIpwRO8QsmN/98wYuKptZrgoOfHxCB3XgjURrzl
5kwFe6wplvzFMsYIQK0n2DLSP4nU6Io9ac31LvT01jd0Y+wT6P3nsyZGVho6njU6
0l1VWa1J14vMUQ/6Gwe7UwpY3VP/0nV1adQMZDxpwL/bz7AWnueLOvFEpwKxTS8G
NnewQnFcOz1+kYpxIVQ5vb22/qro7XRN2CzpVcsyK1+h4HWJPvczDOd/pKaktpJi
dV9fbmxLdlhrD5VvHCfCxAjLd03YOs3hhBeH1bfw2HoLd78dsRYib2HxYwxomkXz
9M8X0lOhmWX9wVDZv/+JEO+4eT0sHc10HNO5W2wgFeNwWgB+NY5N0aejRtOx4X6C
7+B9GavkAZdIQUZLjdoIJNi2sw3e1b03JDU5Hc5wzCD96Kzq8NVqCletzp13Nurb
Aj23XnyebT3x0S3CwkAgFtMUG8i6kU1+4674Gph75FHfcD7ZAsJEzAxx+HjwgJLZ
/tCVFO9Z4Z0zvqwteihcdQ3bUAuuh/QsM32pJMYJDq4V02+yMZBJhKUgjpvlN8JO
e2rDTD90q8dS5JLTUBF8lQBPafbJc7t0ZuziOHCkPBbhQ1ZOUX8l7ODfzty8h7ul
tE3HfNW1vcdwn2X2kKoKVzF765mJ2pt11ldmKgP2nFOpkqFS/ns26A5L0NCYLH2y
05yq9AMQUQns+U5QwgFTEJ/2sB/H5oVCS/xIgobvsRUiXtUR7SAh3lpYJiKYd+fS
N+AyOz2SY3vmOnzCGBryMKG+Jgg8ube3bZgWdvLudzUu2ZFrXLw/jg2ZSJP2UJXb
vvR/z+dLXP9K3mTvsDvdBB2w9O8B05bJtXXp1CGLKWbwwWWtfqAsjikAFeXEEbF2
DTJR0VwibHe/AzFg6ZeY8+ntFbEoQnmjkEM2xz2M32XR2GPDItxUiVSA/Nk8aB6C
+mMhzkajUZncwixKh4GlVdvJ4iU8L/6MkYl7J5bu8PrXrWjwLQe3KrmyVVA+ax+a
DuTTkmSfSxG8FbTi9JNonBwvG60SzXeQTFUP9Xg2nhqh8O7NFUYliE4kpPdN0l9N
lZSBEnQdfeR8hzGq/1S2gDq4Thm0L9zdiO3FS/BPTeQJz1/Uk4o63o+5/Vm/qLnQ
YURl+3Qla6/e9iFOrSb1jbdpme16jBCXg6YfGcwiDJNQdGJxZ2bqDj+D2Bj6RrIv
EUOkfuRpcAGxORV33ayN5dUmEx5lK2PTF1wyhBFlnPBpXeLvW5vjoWhy0gphbL9N
8I3MD1ygXGyfVg5zcnSlXLTHgiRHIeLVr2RX2DDN2XTuGzDUkgeADjLdZhdferZP
tm3OdMXMLwlEPuW7AcLhyriswFU1qG2t95Mo1M/OAbELLpADqw/t7pBeBs8UeB03
gjaTxwVRfYfEBrXcjnnnqmpuwyhnSZBqTTnfL3PrBZrCvFzZRqc6zq1eOmOXkicq
nBlcXarYHnbJatzT8TMoNPoTxbcVyR/j4P0QahfSfgQuJv9TJ4TVB7xkh5+sDOn+
vQF6bPkd2K1Yww/vNNem20Ug+UZuyH6UVGbYaRIUU0FYTOtsJEExB8aF9z7FjZHV
LcS7rrtAUgpkVCwWHFOUxA1jKNs1ZM/N6opfviMTIKwe7Ckk527EJWxQDkL3+dx5
h2YsrSJQ6Tw1DeMFR157juyppljMu7YchCdbHJs8A80lGdqNh9a0CXb7fVuJGkEu
6mHsVYPI4rvddZ7hKCQ3JeIZO4dPk3KSrcEWRY8XOIvUFc6HhfZmmYwdEKOnY8zq
LO+wEXzi38AACnL6EA/4poxA3ZI4PkwOQM/8iAVQAe993wrZFIEf4C3bHSp4hrr/
4K7Chgdru+xiMGksiS0CRjyYgI8ZwFk2x7m3mAhClCSxRC0IGPkCPMA2foO4egwt
1ldqEv58yKAdeKMvfWrzNie0LbCNHizs7SNh48gKsJ3LP5Kx8vk2xeu9f7sNMjOf
205635IFWm0OHJDKQBZJ7TPiGk18W+fKxasmE3lvP4prAnWugm1kHNFxDo9Ni948
QIAbFGW9ps8e2nTk2H3Ao6dqULIhCT5k7M3F5Lf1U7MlI7ePTQALGhOTJTKblW9s
++Z0KNjrvpAVjxnqhtfqeKOp+NBuR8YlGu5i2uw1G0ZvLdr9JcJ9XGRFiZeo7XQo
45LB9zL5FyyaRc+JTMjBtDlJ0kll+3Y4JX65xvCZ1f8dV4f0r6USiQuRIOKMSnD+
eVs/iRBFdX8mfT76TRabbmIea3wcDNNLgRj1pjKSlNWHSxt+ePSe64jQOo0Cm6QB
/nJPXJGutYJlhamhv3Vsa2aHOdttGuz6r4iMTpgR26SsTV7+nDCFucfNNpTZrq6A
329ArrRRPPR9omde1viDWWfv84ZjOP3AnN/JlfGTmacziLO41OHl+EZ9UZOdDYI9
xB/wbTUsosEY7Ad/JUVpOTR8e+VstruuLU2+Iyvan0Ciw4LIbbwIP6UgwXGl7wBv
K03xBq5ysAAOChC6WO9cR+AFYKte6rVj6tDwtEUY3tG7ubLaj3LDlXsIHXsfvMlB
usK56eq70z9Z+L60QnyWCeip4VtZaEL3BJKUMizmc6iJocT0LECMBaPewQYFldsS
MpGjrK6FKLWrrffTSS6nf9BGXcLbsrwcn3JsBim4Dxg95zwykDEV/OG2R72NTjHq
CaUvM1hlC4shjXVIJ7OJHe2GDgr42d22C6q3jD0Gfsk8ncvBMnpg/USdPpmJ8W+W
vFRqbL0okuXCZaGNTWqU9AM5+Cvx1LG/hVlSWz6wO64Kzafi2Kib3ABq2zWe8w34
WDGNnSVnd7OIigMciYzAv0RHyHsCObwgR+Dn3n3IqyDrW/DQdSmSVk8qbrui5bSP
WwF2XM7+1C9CVNm85Kv0AMLfaVmnU2SdjcOrMH4fgE+GQEhvZXtepyP8H8wOpx9O
T7SsrKz0MySv1exmrpltGhyK/YU1zy8YkzegtelBe2eGBcO0zgUh31n4MMlIMWjr
S9SM2CDi1sHwTtobyRK79xzv0KY+RAhcAplFPrXumv6k1ryAe+j2GEdTVvw4U8fQ
T06CGctIzzA4M1RpE/ZCzMYgUCR0ewe5cF+ZT+2AK4LI8h1d8A9wFRSDQ+Cyw1p0
SdX97h3znyKhsqpqGsSadoLaIF4qj+saeYyV29YZIryCmR8Ez1O8zaKNsSnXFi7/
H7hnkXiUGg69mdMJuOeZCEN16AeHagRtkaxoUHXAdD42cTX3IYeIU/BNnPXXtt/e
yPMwzJ9esxDcLue8w5ZM4nRj/s1P6RDH3IyFxkY/uLIe7xSLcYjv5pdpedILFnFp
lLPkYCnpFpFSYwLtQ61DqP667Akb5cCPPjzAZt/bVpGAlBawl9usqh2BUnI7PN+e
Rn4h9z0g4+v2ZUY3mxoLE0UOyq9AgYyxadV5vQknOaaGdvyzATtNzObjFBuvBV7K
sDpberMIYrDsqJ/SeNBoGNEduI0lzBtW/F7HBDg3+0rg2HYy7bHFTJoGBfGMYlET
n4hsDyxmdGk5qOhlFyWAw/udK+N4qaBE3WSTM78H8uSBEZnQ/KYIZfjiBsQ1CcKv
ITH9XlzQNV8e92o8gk1x7PKBIg2Ispz6k6FQIyU1rVaB5Lx8z23Ut1UZ/MuVpDDL
WMc1TsqdGqafKjz0bPsRL3D6PIBVDD3UahOHEw4WMqBEk+li+2fhxA/sBRzwfjJ5
pdv+PrF+vwf0tasY/j6klx3dOzrQPcwdzeMv99FrcubXFepUDrJ2VP+z1j3SMLdv
F2JJndpSyExsRK8ZGPBQmKC6J3B9LWD9CAdmcP6oZ0Wj3wyc2ljBn7L0mp2NdWzZ
7T4O87XMvVAVHayVJLmUVytyETD2NWLPIScEbSY+je9Mrtf3Rhrt9Eat/OfMqFle
9fvA460ZnSOYuaUJUYLNekp6y7JqJ7uckFcjrItlhkOCtFS76vYRciK1pGrugFib
xN+VoGeU5piQnX//D9V6L7Pp7Ci49bLNYskT7vc4dt5B/gzuDYjfQiFpA85MMJwP
7OoXquNzJvsV0d9oQrEHJ9yL2XOL7KaSW+ae7BJasFAlqCnmjPCwFqjdYBL2awCw
4P8XzraMI9EtTUtHkrdL69Y6s7pwYXdm/7aRedRsflq3eLXGKoQWWnp7jCV8oZfc
9TKN2fS9DcJvz6nhyBIo/EqpNNNckQLukGvkBDtRsTcsuzt48PtEIP50nvo3h6cv
0PmSpyKshf9ryL6XT/BYd69+YZcr502QUMjaCrozTEzksYe4TOvcNe8jZZIXS0ki
0uS7PffSeX1zqF8nn/swo59yzmVbaIR68z/ipmRrSOkq1vFYCdeN8l0q7iHoNCRT
pivfXsptAKaWerM8k+IzO0+exyc3oRFumE9CGnPE4b1I46lCUfV3pwvQbiZESYNC
7y8w4fA+z4wrabvGzj6ftakbMaL6eEtu4fKlmbXcEXpKDSihkrYGSRwK/tH5U+ms
YTlmUTPXZTSNn8aZHHPcg4xL9hTMTJ3PchI4CzTn0v+mq773wSDvlmyXkb1BLshq
Fn87MAiyP/7IVnW2jNHst4ZFNKDinhh+OHrkV38nxzk7EJwqE6cKRHP+LX3Dyi3n
+k7jv7WeE3nzZrx0V6Aw1VZr9Q8uohcByKFL8RtzqK7h/he+AqDlChCPKbqHhKdN
1G4e/5Gl18tNH4Q7yFZhddll4skRu8G4tdA6hREYifnuMJMhdtvFslIrF2bAPLg1
gGgv7lugPn0etkd/CLTHAepe4o7INrSB84j7nK6H2nblKTb2tzzKntgMzl6MLHWd
VO+owLrsR/R6rMuUtzSAB5r5B177ateb0MYxWggt+Usj4tRgwXj2yZrDVMtA4D2+
gR5O5t0L5Cy9lNF6R8txvPW77LTTas19TJxt8lwKNnGQnfdWVmWuNJsACXxuTVdA
ohU9l/cHw0JhYpmdfJ566VxQHo6iUTbzRihLQQgwp4y+penK7kaYCXWkWRxruURc
/7VISuNfm9VbG+TI8mxKmYUXHADFxvwOtZ30q4FOS6MJiTb+wBS5Tg1wHbieJG2m
jQUiBHmge/rKgJhhReOIATbzYrcR86UnTatvDEjVYypYXMleJWlI0TDanwnBAblV
YUr2DnjpNmDzTX9vjhEVnLkoVDqGOvbCJZxdTK4Q5TGaPV9DlRQ5r4WqiwAYQ5Pw
1RcIFH05YDiki9BmECa7jzCvCKQ5ag1w0Zha9v1Ak2k2ieTdD3P3tXa++n910Jty
Nj1DlX8zGrvPfsnjfOAoQblizCCVE7xhq54uNhbgLk208kC8DHFCLQMFL9x4/7cH
BBemAqbGMKB6/Q6K2PT7zxqIXN8TLN0dJOaFdVp9Oak7ydn1O4ZRA2d7aDrSpa4M
uJI3XqpAQzoqQ/m8WLaGda4dQs8D9Ftwh/6X4fwJnxmk8vNPvKl8C6hPiCy3lXCR
SDh/j6f8LHGjrnTtwwGjyYfWo61oElHCrY3vZctZg8LlwtALIgNZJgh4RTTBvn0D
01HlHNT4pRqTY1ARLGfN893ILgqFLfkJ6Ie9auTCAheZDQQsSLW/AZpPNOHhumSS
KQZJz3CAHrezEvwe0k5JXneQNYVdBcDJr2pDICJjK2M/i8Bzngx4wVTbcKMciWBu
ung7ZAIm7Y4MLmSY1+tdfol+T0y9VIP2zgqgc4E4OjVQ1HhkMqtFVuoyvUHWxTyq
zRd+G0eILgEmjUo/WAvaRsNeqeljqiHgektiWo0IQ7GVUh43j2B7tStyWp/YH0P8
PnbmRtktV8fLNqTLBiwHRLxudBFb/LDaaWd4WtmmArYBfGFsgrneQcM6XfoOgEKR
ABcmfFgIzQvvLPN+jpDeYxYd0vd5jJNVqZg9wXRefcQ=
`pragma protect end_protected
endmodule
