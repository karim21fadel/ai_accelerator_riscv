//*******************************************************************       //
//IMPORTANT NOTICE                                                          //
//================                                                          //
//Copyright Mentor Graphics Corporation 1996 - 1999.  All rights reserved.  //
//This file and associated deliverables are the trade secrets,              //
//confidential information and copyrighted works of Mentor Graphics         //
//Corporation and its licensors and are subject to your license agreement   //
//with Mentor Graphics Corporation.                                         //
//                                                                          //
//Use of these deliverables for the purpose of making silicon from an IC    //
//design is limited to the terms and conditions of your license agreement   //
//with Mentor Graphics If you have further questions please contact Mentor  //
//Graphics Customer Support.                                                //
//                                                                          //
//This Mentor Graphics core (mcan2 v2005.020) was extracted on              //
//workstation hostid 838626cb Inventra                                      //
// Copyright Mentor Graphics Corporation and Licensors 2001.
//
// m3s009fg.v
// Address Decode, Register file and Output Data
//
// This module shines out register values through large central mux
// Revision history
//
// $Log: m3s009fg.v,v $
// Revision 1.13  2005/01/21
// Clean synthesis warnings
//
// Revision 1.12  2005/01/17
// ECN02374 RTL lint warning fix
//
// Revision 1.11  2003/07/30
// ECN01958
//
// Revision 1.10  2003/07/30
// ECN01953: VN-CHeck code issues
//
// Revision 1.9  2001/09/25
// Unused signals/registers removed.
//
// Revision 1.8  2001/09/25
// Tidying RTL files for review.
//
// Revision 1.7  2001/08/09
// Changed 'sl_rx_fifo' signal generation
//
// Revision 1.6  2001/06/28
// removed unused signals
//
// Revision 1.5  2001/06/26
// Change sm_exit reg to posedge
// Change state and associated signals to 6 bits
//
// Revision 1.4  2001/06/21
// 'mod' re-named 'mode'
//
// Revision 1.3  2001/06/15
// Register sm_exit on negedge
//
// Revision 1.2  2001/06/14
// Files tidied up
//
// Revision 1.1  2001/06/14
// New files
//
//
// V1.0 - synchronous interface
//
// Include MCAN2 states
`include "mcan2_state.v"
module m3s009fg (xtal1, xtal1_in, wdata, address, rdata, txdata, rxdata, nrst, val, rd,
//*******************************************************************       //
//IMPORTANT NOTICE                                                          //
//================                                                          //
//Copyright Mentor Graphics Corporation 1996 - 1999.  All rights reserved.  //
//This file and associated deliverables are the trade secrets,              //
//confidential information and copyrighted works of Mentor Graphics         //
//Corporation and its licensors and are subject to your license agreement   //
//with Mentor Graphics Corporation.                                         //
//                                                                          //
//Use of these deliverables for the purpose of making silicon from an IC    //
//design is limited to the terms and conditions of your license agreement   //
//with Mentor Graphics If you have further questions please contact Mentor  //
//Graphics Customer Support.                                                //
//                                                                          //
//This Mentor Graphics core (mcan2 v2005.020) was extracted on              //
//workstation hostid 838626cb Inventra                                      //
                 cdr, btr0, btr1, status, cmr, mode, tx_control, monitor_can_bus,
                 ocr, clear_tr, ier, ir, txerr, rxerr, ecc, ewlr, arbit_lost, arbit_lost_position,
                 rmc, rbsa, acr0, acr1, acr2, acr3, amr0, amr1, amr2, amr3,
                 bus_off_reset, sm_exit, wakeup_int_en, state, illegal_sm_set,
                 sl_rxerr, sl_txerr, sl_btr, sl_rbsa, sl_rx_fifo, rx_fifo_address, addr
                );
input        xtal1;                   // main system clock - ungated version, xtal1_in is gated version
input        xtal1_in;                // xtal1_in is gated version of xtal1 (turned off in 'Sleep-Mode')
input        val;
input        rd;
input        nrst;
input        wakeup_int_en;           // wake up signal from powerdown module to reset SM bit
input        bus_off_reset;           // device is bus off so put into reset mode
input        monitor_can_bus;         // check when device has begun transmitting
input        clear_tr;                // clear transmission request
input        arbit_lost;              // flag to show arbitration has been lost by transmitter
input  [2:0] tx_control;              // transmission control bits for state machine
input  [4:0] arbit_lost_position;     // bit position where arbitration was lost
input  [5:0] state;                   // internal state of device
input  [3:0] cdr;                     // clock divider register contents
input  [7:0] btr0;                    // bus timing register 0
input  [7:0] btr1;                    // bus timing register 1
input  [7:0] status;                  // status register
input  [7:0] wdata;                   // input data
input  [7:0] address;                 // address
input  [7:0] txdata;                  // data from the tx buffer registers
input  [7:0] rxdata;                  // data from rx buffer registers
input  [7:0] ir;                      // interrupt register
input  [7:0] txerr;                   // tx error count
input  [7:0] rxerr;                   // rx error count
input  [7:0] ecc;                     // error code capture contents
input  [7:0] rmc;                     // rx message counter
input  [5:0] rbsa;                    //rx buffer start address register
output       sm_exit;                 // update reg clocked by gated clock when clock disabled
output       illegal_sm_set;          //fire interrupt
output       sl_rxerr;                // NWR strobe signal for RXERR register
output       sl_txerr;                // NWR strobe signal for TXERR register
output       sl_btr;                  // NWR strobe signal for BTR registers
output       sl_rbsa;                 // NWR strobe signal for RBSA register
output       sl_rx_fifo;              // NWR strobe for rx-fifo
output [7:0] rdata;                   // register contents from read back
output [4:0] cmr;                     // command register
output [4:0] mode;                    // mode register
output [7:0] ocr;                     // ocr register
output [7:0] ier;                     // interrupt enable register
output [7:0] ewlr;                    // error warning limit register
output [5:0] rx_fifo_address;         // internal fifo address for CPU write
output [7:0] addr ;                   // feed around wrapped address to other modules
output [7:0] acr0;                    // acceptance filters
output [7:0] acr1;                    // acceptance filters
output [7:0] acr2;                    // acceptance filters
output [7:0] acr3;                    // acceptance filters
output [7:0] amr0;                    // acceptance filters
output [7:0] amr1;                    // acceptance filters
output [7:0] amr2;                    // acceptance filters
output [7:0] amr3;                    // acceptance filters
wire [4:0]   cmr;
wire [4:0]   mode;
reg          sm_exit;
reg          srr;                     // CMR bits
reg          cdo;                     // CMR bits
reg          rrb;                     // CMR bits
reg          at;                      // CMR bits
reg          tr;                      // CMR bits
reg          sm;                      // mode register bits
reg          stm;                     // mode register bits
reg          afm;                     // mode register bits
reg          lom;                     // mode register bits
reg          rm;                      // mode register bits
reg          can_goto_sleep;          // flag to show SM bit can be set
reg          illegal_sm_set;          // illegal setting of SM bit
reg          abort_transmission;      // upon transmission error dont try to re-send
reg          single_shot;             // only transmit message once - don't re-try in event of error or lose arbitration
reg          set_re_transmission_off; // disable further transmissions if error occurred
reg          sl_rx_fifo;              // decoded write strobe for rx-fifo CPU write
reg          sl_mod;
reg          sl_cmr;
reg          sl_txerr;
reg          sl_rxerr;
reg          sl_btr;
reg          sl_ocr;                  // decoded write signals
reg          sl_ier;                  // decoded write signals
reg          sl_ewlr;                 // decoded write signals
reg          sl_acr0;                 // decoded write signals
reg          sl_acr1;                 // decoded write signals
reg          sl_acr2;                 // decoded write signals
reg          sl_acr3;                 // decoded write signals
reg          sl_amr0;                 // decoded write signals
reg          sl_amr1;                 // decoded write signals
reg          sl_amr2;                 // decoded write signals
reg          sl_amr3;                 // decoded write signals
reg          sl_rbsa;
reg          wrcyc;                   // read strobe
reg          rdcyc;                   // write strobe
reg [5:0]    rx_fifo_address;         // internal rx fifo address (0 -> 63)
reg [7:0]    ocr;                     // output control register
reg [7:0]    rdata;
reg [7:0]    acr0;                    // acceptance filters
reg [7:0]    acr1;                    // acceptance filters
reg [7:0]    acr2;                    // acceptance filters
reg [7:0]    acr3;                    // acceptance filters
reg [7:0]    amr0;                    // acceptance filters
reg [7:0]    amr1;                    // acceptance filters
reg [7:0]    amr2;                    // acceptance filters
reg [7:0]    amr3;                    // acceptance filters
reg [7:0]    addr;                    // externally latched address with ALE
reg [7:0]    dai;                     // Partial read data decode
reg [7:0]    ier;                     // interrupt enable register
reg [7:0]    ewlr ;                   // error warning limit register
reg [7:0]    alc;                     // arbitration lost capture register
`pragma protect begin_protected
`pragma protect author = "MED"
`pragma protect author_info = "VirtuaLAB"
`pragma protect encrypt_agent = "RTLC VELOCE", encrypt_agent_info = "1.5"
`pragma protect key_keyowner = "Mentor Graphics Corporation"
`pragma protect key_keyname =  "MGC-VERIF-SIM-RSA-1"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype =  "base64")
`pragma protect key_block
otlNgNcv1RJyXavdJRR6pM1v8TmIkSQnJ8p4tGi6lxcU9mUqHm2yIwPK/CNHU9E/
dBodbtP3k/tJK9VTWuLjcwjW3diKZPlYc8uPdVdgEmoZ2elRXLj28R3tl/vR3f4m
Pa5ZWm4Qiyeav4/FBAt8CF6Ab1jImptZyJePF8kMRGc=
`pragma protect key_keyowner = "Mentor Graphics Corporation"
`pragma protect key_keyname =  "MGC-VELOCE-RSA"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype =  "base64")
`pragma protect key_block
qlk40b84zKqkNpYGAmpui/1s6djMLm5Wyq09RmLJRo8verh3kDWDk4ukcpsr6Qw4
ESP2Kdnctk18mQDwYHST3+b9Cnb76wP36RWa7lYTZwtj8QnOuXMGUfAetSo26Hc9
0O9ANlqHP5Lck9bO83bAG/I/psTQL2gdDns8wF49gpA=
`pragma protect data_method =  "aes128-cbc"
`pragma protect encoding = ( enctype =  "base64" )
`pragma protect data_block
IUigHciSrh2w9s+qyBTAmiHRODgzw33qCe1YTeSh2tZAuvyl8cctX5JmZuFakz/V
4MRNfQTJRuKC3hcWaMUfQDqmTWN08Uo2jyUSftFKlhuO6146MkhQlo1iocdGLiyk
4ro49pSkzaah2zXyVGXIv7Aytgi3b+JvkPfbIkagZSmmwYuLN2mqZ8AGgOx/RTE2
TGjuntyNGr7lH+eqRhxj0+3TJ2H1GE1xzgjoPdKZZfKQJBmmxeIHKNxX5VnCLXuk
1Bk0ZjlLecfjO7n3eDyStIuDhMahorbxvAEOig8WvMGPibd9LrzpKXaLPEmneRPv
c9Y30YcbrlTtB86RsrFYO5waRxyJyGWntxwe0VEcQhIWY0/4Oj9jYL39I8BSmQLe
ENsezwCYhI87X6Io7iSfc5dHwu/h3dVIk5+aI0+mSwDuxvGTDSMQg9zeNM/YkHNI
/WdBdXmi7mYPVJ9cQzEFIWbN85yVzpu8Pqqlsyx9dTSqT8zyW84VT1dL4md668pt
xij1SiIBkOfWa3lGmI25zdlJZ59dVFJCXRAd5PoQKhney47pBfj5lyp+27/WBO6Z
bRhIQ12wS/5WWmNkBLq8pYJkaHX0P7LbLIsukWEtPg/wFN1qnzHQ/4rXv6GYhyWF
36YSnPOeTElWxOyAZat7CAqRHgGSzk1UZXUhTdx31soyYBAatjerFiUGqy9slBph
nyKtVDxnHnx5nBrHhqpG7TudlLaycqH8I7MGA88hr0BP/wOjUZd3opX6ObEKiBrO
5pMnC7XndewU6OLAVh/FlVHefj1F/4eT8qVX2nOz2GUO7o1MEDTVN/UGrxOIR3uX
VEGxayDJjGeUIIelfiP0UwPt62/lgYtQ/HPLsR+CeGYGikdO03ZYoDHaiP5wM1RT
3Q+Iy6+2o2pICqkifn2zN40EsdKDAIA8dhJHISxPPx0NmRA7n9YXugatCS1DC7gw
juur7SvP+OuNNtWPb0I3h0vqQExmGWZcCLx41FqNj8a/zndMbAY3288GWtpnl47d
Qq6g5CG0WvaLAg7vMiW7d2kU2G2sbXHM5/Go1m2yMjNECGLwWf3crBytnSYO3WDc
H/GD8E5l7EA8FencBEefUEEOm2z84dsZFl7vHOnuQ0zymkO2/8A1WdjULq8vyVZa
OX55qX8HOfsd59Egu//Y+X/I92HOcapwRTHYz2nev0hH8NUc0Qf8LXI6vYdZUMss
EbsdXgSElARpP81y5OKwYar9KYFEockFjd74/HD1k59WeoBK1CFmMlNGaOmrVXhs
Fdlys9aVX17wVdbvrqg4ktfWv+vLAfk1hTYtZPFitgQPRX15SvMt3jNHUMCeLpme
5Ao4objqrMorGszXrg8Dfdhn/SxSXVfqHEMXGoVeOEwBgt0xjSsW3SAV7lypJiEx
cm7hkAJnLYRwzkUvMVTlJCm9a9/EpD2la2IvEaaqszasRod0FaqG37ECyRIoZVUm
ACIxJ4rponOgvW3cg9wduSUv9zgTa9mBomsVa3RvrvZfGndBRSE828a6+rXXTbPo
nLCkY6psM+25Spala1WiqfoHxL5g+fjdlkCatQM49jtj3j+L0DGTtIYRCsH64eyH
et+ZB9Uyd+G7gOW6F9V2l8XmKoGjQ7Kf/FAC2bMSIABZySi2EkLsFydWEZeabvpm
LPxTF3FFlg4F01m1J27nF/1hhT8r+ubfnBs6IqUMmVUcAKC84DVEkrfhPZMx7R7K
kxioKenCKgnw5VwitEpqOwwbN7KdepOebkqXgYlYikLvE1Zgw9Km4yRc3lOnufHi
9yrsCPynJL+WOfS+xZoazSowjmmVpBbNn2HOvr3eLhQ72SWO7YjilGxhARk6kHq0
mVIVdcLicVTXUg75094xm0p6PT14TYX4E9dxhDHJcIf+sD4gK6DwF2Ogm07zOmQS
xV7IUfBiCwJYSsSMiB1YWNpV9NtrqlXwyi7cuRyZyxbdREDlGYns6fsJr6sfWZ89
Dti4q9A2zg1irNdChvKH9WmPdG0WCEFGKbm4SLoirRCZQtYtadS6TVtSB7IQwKUN
Y1bjuqDAF/FqOiMOJjOHx6ogf9rIYRlrxzQoLhbaNjQDJXeFwqTqevfOhYx8Jbqf
uJhARzheeYUtGl/QwI8Ovm0UhGi6EozwWdHLuuI7oZfEJwQC8I+zg7kiRAmg5dI5
6ndKbW+55J1OHJa7/HtbaYKEF/9kyOstwj9vBywZt07QUkXJn0HK1V7v4BUYRVt9
++T2K1xFi9uKgV3H4O2XPMHXNrBl3GRmbi+/lGByv5NPso67tkAVp/s5KMZNHxIZ
dVHtR9rgQAnEiJdbnvkhu++DlSAzVx7TiolisJY7jk83zhCiw+SonLr6Z/XYekb9
pYQdy+reBkDAvAD+bkzTBIQrx5JsEUvVbaUVxjEm/tsZldMFDm+KP5igIZTzAsOs
P1t3k4UQqLcIu6OhiAk+9dx4iXJNykpyBFYgn8B/T/lE86pb3wfJKmdfHV2STDli
/Mt3JZOCh0m3MwPE44Opezo7e0ZKurw/0PtXN8NLkWVoDzTYTA9ftxyHSjDG0g70
hvTauRm0VNW0jkdmVACrsr5mOdImlZyteDt+y0vgTDWDl+ObIPzokIxuFEk+FKIp
0ZIi+WvnAwsB/YRBZ79g1Gs54DrrC0pr2rSmg7DgHEnO84yCJIcci1LZN7LFwVvR
IJa4/T6wYYaa+Z3wh92KLdO0nHUTPxyyfjwu4Iom+2pV8HkBKVWlmIztDpcWti08
aN8vxCrdrF7Z3ZbPmjMPSKpl5L9mtZYLe6a1OnLvatrU2bipfA7MY4wpdPvkbF6L
QC9wk9OyD+q9VYsVcTp18EqfMFJ1rg5DlDZUkLk0xeLXvlRquYON/EbjOn8UEu8/
dAc1FTxj4r09nU4gtlyJ679fuGQ7JLEWGO1wke3VC0oSXYPJchhsoT8cjc/Ct6Ns
T8ht6XZKevJ2PCHkt38ch3F3hoq46NXcHFspO4pvSMB0jhR6laEeeIaOHnXWeOX3
pnqtv183JBnupPYCm4Szm7CtPGoLh0Bay/uBm6VwqTkr61aG9IelOkScYQOUuOIb
sE9LntDrQ5yqOrE0Kel995EyEzRsNa/sLTcsn/ZlfaGj2cYXG4Z9ev08cngDXZH0
n/fsN9HBPp+WqzAKRGKU60Gnr2kTXPa3SL5GohnvHJC+KNRGgJXiWOse29aKrtUM
ShnI9pqr7EQXEXAR305GT/NiO5icntAt3gPM8TnPuRZAt9P4KQcQGgXBHBkPVKhl
vNWjHBriKojA0qwF2kOwBYr1+BA45Fj6geyuYnP/9yuOjQAsFiY+FW636cSUPugb
ajS+V0vI9+ygSzfc5vGiFXfjGhxXo+48lNn0un1ohTyoMxgPOIHzP054KyuZ9zx2
cqVObttzNbOjU2Vjev60cD9Wfl+VKDW2uqZWGX2ZaaFW08knA+9GfLnD16+smvdk
T/Dg/fSgZ+C2MI2qdazyb2rR9U/YTDPiFfPRQw8XJJET7eIG65Ws5sA1pFwCfxL0
pd324z9YUZqrJqrsbJB4HNapGJ5X+OXokNI2b8wInYaBYYlNJWCzY9WX4n/0FsSz
AQTvTIOOHekxwPhNFgt7/NlmP/hL0frQc4p4ahbDobqe0ZqNx4C9y7ApzUP0fdie
s5L0L3rMN2zxa8X6VIlPBA6cKEe/sLJbsBURMIDMX2kzQTWj1238Z1pLeGjppa8E
QiuduvWjtt7QG4eTjN4XVM//vELzDDlcBqXk8wc7t0fx2YYcmr7bBjvwN+4PHEE7
DuOs6PMlEmFaWNMLazFcco7HIJ+qi6J51cpXnamj0ge3k7EQwbRsnb/TaWHJEFhr
AM6q6P4E8ov4uGWZrsixn8VnyAEcF6kUXW0J3hMUSBxMyYzykH13cnQmijy9s7FR
bg29YXilzGlrWxpedyxVbaqdHUuZB0uE7Ln8dwQEgX30tp/LaEj86b9yRJo0vUSm
5KR2gngwoo5H951S55mahvqqcnRZtzFnZ3x1YaiVC7CGNz0eAsr+iRkwFoGjdV5Y
aISyqHEG98q+qvImKET1KlJ3V+s4J3WaVpS2ulmzjjUig4zoz+lsYvuHt2AfMMrv
Eo+SHo/aRFWZC76oPbUFIHKwIi3LQv+FCzmhN18ev1rLR0amv7SYqD9bO0M65AgM
iaTwyz1oyDbvLYPqzt929adNAUN85mQ4PecLDLX9bEwfhcL+I4Hf5ROTnNSSSj6k
8p68iKyY+ySqNsKjF+Gqe7zUljCRcRupHhmq5oLLZz3vEHgFgutVphN2Sy9hEugJ
BBnr5YWy14fLUmvEfyCPFYGZZ4/MCQd0W7ThH+eMZG85AI5yG8xnjor5nPtF5e4o
JNdTHeOqujkWHzqCBnjUTSqKTaApReeQgHQgGWX4XrZjzo1cYOJovyqTNdqT18wE
xcNGysf5fg8hQMLStXxuWzyLNTIw7LaxuLqmhpLGzikq4yDK6d96dK/sXgheRede
A6UpMX7kuY1MLXVDrzo7ks8MCifVnVynCtFx7HLwoijwpGzIRXpFxBdOKhzfXg/e
2SgfBfFBv82EW6lWDyxQAzza9w5jafzTo2J0+B0Vt7FDRBzXKXOe5AmI22C/4057
IjIq2lN8mueO/gPsBm3VlyUx/BPZ0ZsXfb4g/hvscDRIt5x/1s7akfKXKb3+h8D1
sB4wN4p/xF46ztBeD1Qpbt2tK+TNviNkmTuouK8NeLHCkv7ut3qMupO8FXUNZuNW
NCg4cegrlYc7mbNqfHoZSphJ3SS0br9QAL3VrH16UQsm5+updn+NP++sCyLmhScm
hUAxuZ4ilnLkZZ3E0hCRSeEMF8lvgK2xrzMN2WeEcQg5h99jn0X5ffAk6RKGSql7
/+kH4yhko+2YtAwwQyn4B3E/qMV8r0OD4LyGnUzoNY1XpUYrxDLV6U5v9olRE3i8
a86myqJaTiQ/UpNZBSBvrcp6QyGGH9bb/WxAE1XzpJzTP/Z56FFrK/fqkk90YLp0
6IL1eWAfJtS1C93/V99aNWengjTA0i9QDe8y8eCjq0w1FWqmRKp0AP9HGH3+P3OB
KVKsnAgiJ+6e2hwp4m5GOdanC2k0NjjgTQyJ7HV5IHKOcBa6+2LHsQzEPsuSsMNv
QrUxdlXMEqgn6EnYYHKhrWsMx78HbP9iTPQMlR+3ifAD5ebRmyNnOHQvgSYajruy
Z5pxLFTWof0BWAlF7fK6mxOuqqR2lFZs2rMKbR8QKtla3H5Hf8rymtonp5BDEuut
iquWmk9fsZGdz3X02ndMkgNqpyt5LLkdNYqr8nDXYsjkg2rNEB4XeaEg2yGHaqWE
8wzLmFvkb4qMPHCRhD9LZQmrQSRtkOPELy8kTVzt7PBK6RAX18whaYSKXyXdSkFw
XmsMDGcmIaZFrBcJ/GQ9sbyFdPp+CV431ILi644McaXM7daTdr+XSvwhB8VBmFo4
V7Ks+xMJ8i21VQ/f3XvUTaISyJSPtWqaGhd++vrhONiDRV3W1kWAx+Dz9wLJwPiK
iWcgsOcy/2mdXNrDcAqJURVYa50ZVhUAWscJDrcmqR4h7dFx8xG/7wDf4yFCKvbx
dSnvwQuYjEkkcmHK8vs4lJhA2vnh2FJy3Xn/ib85nMwFLPq+cV+N3Ud2GSdMvL3m
DarmOQgpIL3Lmp/ARatD4B+BiPA/5LUj8aq5z4Q26LBIukcNpyavF0dMBUosVpvy
LQy719nAx6VOW6X1ldDgFF5Z9TTBsVDCUSh9SruQI4ibkQC6KFTO/0+1Nyc33L7p
8OirKuigCALQcvG88NGHb+aDkPmXvjOyj4zWY5JZPi0UcuIYaDuXbDhOWm5rts2N
8eHRMYiQWNGRf+HSUqE+t9xq+zBmuWX0gVScRDDX09VBofhU3vXsSQSHiDVOlJsb
C5OTXNQfOzTpaqF2XiMgPB3A9B46rl51aH85JyzTfQU8Sxet7hbdcIHdoEGxVCqM
s+QqGqNUBYQyt2Bzhk/JDkmdV7enxMVyQlopW7Q0zKY9Fng5wW7F2iZg4d5Q5be/
AV6sBOGXQ95w/kq1Zrr7w/OIPnfgoqO/T1Mqr9e+d+ylt4WbQ2I1R1We1pmsuKRz
jBSpt8ves4F0+l8ubS9HvuRu4Xds0ckB80bCQyZ6q31ba7+C2F4UAa++EWRQub7g
rA3rm283nXFj7K0Nl5Awyrdq1dsDTIa964IIgIugdkg70c8dYm/wY8fpO6ujfH9H
4xnZh50IGKKXxmwlu9kN3JKedTOPGtEbC7ah+PJr7qe4fsF3wJtpeSVRIbrtdmCC
dZ8immNOGlFi+PTFpe9u46njWXYr/wC0sHrJx9NPf4MhIIpIQgND5zdAyM0MlDJh
frZ+4/KDye10o0nWKXhKHLBdg+vAcSOBJmcr9ja5YQqGfE41FbvAJGJQtSJroIq4
5l5YveJQg2268C6mfHaFzLmVC9Z5X3yNPoEuwasmymI8+PWZx3UE0L9ohfO8HD+K
XdSoJ0lbJMPfPZMHn029imc2RqG+STLFXYkv4ThG2awU1FUlQa7GiPm83uMXF+Ah
g5rXnsh9zogOlLggcXvwYWkvyn7TRm+qcYWCNejqVZsxcyZJZzrRD20k/WIQ6xmP
NjUbNisrptZ6TS/QTXp6AlW2n+FbIvX8DnI38+rjK3mcOQIObFGWm9o4vSlCcx2T
/ywg4MLzGf01XhJciBmnwKTA1NIPBzEG6RkRqbHpHI7MQGTb7+F952mk/zFggPkF
qDPqo40faMhiome+4E48DPIX1pVjvfhg67D+J2/U+adTww8cySnh7U+kcZ7mrdFa
qu1gtZaH6TDlo7OawTohl3hnuJb6bamUjBBuKYgCopm67A+NumXGdNt/rGE/8KIB
cQ7xXDbXGQebzukAjzrhYK09uS4E7F2wPbUvUDBq3V2rNyBV0MVi6Swo016OUvXU
n/5c6aVenEGBpJdsMj09C82JDSbL5pRqxRnAn1UlnV8Ru3rFMFO62gl5wk1cq4Hv
IRZdELM6wlO4xQl+1bAEPq0ctY4e7ktFSBEKy03b7P0m+mIVwplxOlR/7AkFlRIY
ENyhGJ3LEJtHy7Vm/0wwegfv/8h0BvdNASYsiiR5RaruVO7ck/5U15az4YHAn8BK
YFGlhocgQ5bTwGSaqKf3H9bJLT3ro3TocYkVupWTNh9TFigFBtGHyKxbaR2N36Cm
SJuDptFYFsKryv0hSWiOysBakPEElFg/uJvkiuwYUj5d1GUNMdl+hDfCs5FGUgr7
G/pbO2UdLS78OLv6OLjax8ufdWskz5RQqtlAVr9EvheDqn3A8hvBEAUSvUZdqpOK
UeMf09Wo4n/b8k1wbxkoWkYtMRryU1v7mwt9fqFdiDLeSs6LuQi+J4PFJ8yj5E+X
NTB9qdbeNbgCc/ucke+yd8vk5D1TYgHWjeUXG8RXgKUil3WOv6Y8D5nyJzS7czmU
2vEYyhSO0UYVK5DE3g0CQVLgbQO/Nnmmu9Dgfgnj8xA5jV+EZ+gG/fPbX4UCXK2q
f+8bPcoozZG03/HC/xG9TTg/M2NtJ4hfSmjklbSBycD2tnSE0w7oeoQJeNVsix8j
dVaPdmUs8Oy5Y7yeWZZAMxDfxF1PTR9jHIecPb9iZbP8soasB/ecj9JXW/QXs4FL
beyQ3VcIrurftsLZqPX1jv10tPmvyaWvPqCbGL+vIdbzB8d885QNXHJOIcUq5oWO
aa/6JuKMYEi6lcvwOSIYIBOMfOO5whclauUOxFyS/QtyQmv7h/YTOAOdkFUcGR6w
U4YQ/EkVGjAGecEVqd7wfrg+nnQooV3SA8ofyJRA3lL+Ak3Z+n6Uk3uT9nGRufX6
+A6eIqOJQpeVJOuPYJQTCuRm+uJjo7QQYSZDDbCxMmveyDmMdJVfvSj3ISgOqPFs
Nh2S93ALaDhG6iMOFb4uPYDBfw/smwKdugJ66fK3D1vD6GwerUV2cIkGLMYTDsBh
JbW+vc4NXRyjv7v0SgVZ07GJBymJQpC8GQAO2a1jvGrOQg2aILoq+SHGumYOCFA5
Q2zpAFF1FPD3ZomSZ64KCgRaZ8+dj0sJTxZmZeacOpidB7+OUkpWsOa06Sd/oZnC
bE+kLqudMenmEgJ8eyIcUGdmfT3tKkMFMOqO0Bsd7jWqi4AmlKBsMJx6yj0HL0sp
Tgj/xYzpqgdPzJW/WcVWGoMR6C1va581exDK6d3zncyCqn5UF5yr/WzdEv0vODS9
CDkZy0v5YRZoeQkYyf9kITPnRDpwofP8039ortHjeH3hcmZipO3qODELHvyx0QAP
AfoO7PYejkTRO1enPfDsUc09tPJlGjzuT9bKy6rR6QXBP3cVvLIYi+qP4byKUTxk
DCyxgY9YIHHE432OUGFgNAdt09WOFgYc1Zr6nMwPV0tOAeeT9NCVQf7ajZpHLp5c
cJzqqz4YrDz9pjVC0LjyRewP6duh3epxQvXG+Oxo3hIoZkc2XyzPMFVREXuE+P+/
nSQzCAzGUOn63dY9Qa/aN3/W7qhF16ZefBEZbWDhP2R05WM78n4/4YUN/8CYv8W+
DrSApGeCYMVZm5BwVK7wWMBdp9m4ivawpjlMvhoFCABfuHZQVnHQexgzGQT7OXdW
YUKbo1rpWRDNG73fgSnUCGNPgOc4I5ui5zvLOUYp8F/oYTLQLu0ckJJVT6pBbFrj
YBM4znb3Iy099cLmEpMVMcrWV1KQ5BkgWsDXJmoF1rgSWm+JCIF6yGuWeAzS+rBH
49Xm+9vMpVU/dj69YA67cvpb/Xp9FT0OSFF4v8Dh1MD0gGorepth69GL2hl1wTw3
R1brU/htyTd8UFmww+dReKzxdgKEl9xKGTnoktJMMMwcj1ebogY3wnI+gfnXDycL
1xaO7w0foUZPzjuTt5d+c+/ARUs9tIHVpoaydkncVc7vz9y6wmSh/0zdaBMY8XAT
fCFXw8Bkzwzlk9HcRaWyQktYhbXRSn6/QRNFaXS2/mQV4KKrQ26HrfycU5KYjhFR
kfB9IhWou1qEr5LieApqkbL7aCv1cWOWH25rkzCuHPaBp9brIDIhN5abrEquCpzK
ltASdsPo/aH+I/WN1EGm/d0Klq26FqRF1QLDzgXhwwhML3XA6nvMD312TMX2G0h3
xniUINCrehrxAuEMS26xUMwIBFt5FxbaiMvX5v9VRr1k/ncey/oudUMqdmAO5xls
7d2shT6v9OvSpL+JgaJOLepto4CnwOYf3tpREpmlRcmKIspoesODraLjjreaM5Dm
EzRYlGgUY7qjXBRCJi9ZhnAfX8C7Dj/8yloRSJt5g9CEFW/WEkEJBju9lh/qW8TX
DVQ/uMfwFzcK6IDQkTwLctFGH0ebuZBMgodXPV7L357KihlIecEPJara4j5a3JyP
qkewuR6Fy42hDvODWtDKWt6ecbbxxsQU/z22+jPz43kiyjPByUykik5eO8m3nDI+
6zdZdhhHYTCuqeiwnTstpYXjvOK2sAM0yudcDNbR+drbKk9k60t48I+OLl7Ugy8a
x0iHJzZ4xlx/tP+XrqcXdSORQOCrLDWWy3rE8bNQy1RmsKRfXkUrDggnOabH8/zC
tmXfxsxuvnyZcaGB2parkOnqSwkJrytW5qUIJMmTaLVZzzCxewI2pVGULdp92nXu
c0+IPI5qoaSQnujIq8JB7K8NNKwaN+yqnZ3S4y9N94OhSDyDSHG0T2jjGblEtUoj
1rGTBQthFcwrRI90FAqkjz36FZCv8ODtn71zk5k6FvGDPqyZM9pdDOtkf1WGwX0g
Mmv8PSx02bb3KIjv2dtOEi1J5YWCbVKQWVDXgHjxRulo6tDqLWOW5K6W1P4dRqfu
9fxQ3Mbs3b4IoyvKnpRkLHHcTjNSHE3KQkoc+b5tHrikmHQbNpxdWRngMNjukPhq
g5Z/aXeyzCpSZfVtzenqONCRip5U2KR1wMXGWMLV/t1WCi3EVHzZ9F1nq2n5SCjS
lXfxgnrDWrvpzNyrhxu8nhCa0l84i0l43Nib6Rh2mru+yrJS2DL6FmjYIbvs9LKU
WRNEVcdJs6RZKMOSRMZwzaF8J8vb1vwnv7/X9TPB37J5N79/J1HLerMR67HkOukU
nYy4WkyQoZlACkyKKcuL00JlkjWX1boH35jPhvB7RNtOr5OhVSLCWn6VK2ABuHeh
xfQIz7Vd53mgApA2UTsDv3SkhJ3YvPg6ciL2rR/2RIj1rfCPaqXsMcYp5qJNt4F8
covVDugsIlX+vb32vwkoasxqj+JXaiVSBkSZG4foLjSzbBiuywNH3qQN5LJ09WFq
xHwb+7tarwYlyyxma6qjKEUqw5KyisjkXXGvIHLoCDqf5RZMXvh6nZEYblAzi4Ac
b0VCHJgqGMDQUKm/7VltrMRAF279FrQApF4cjenlgiuLFDmJlCG33GaSdCDEBSR4
evCrBYYwJaLudqo1Qtata4RhxQdp6K1/17pU1OcEWZvAQ4DQOhdmNaYhifC0tUpU
sW4dmgbszEEer/T6mFC1eOlL4qEl5aSt+K7tvgdZjCQsAweay8haA0CZSqCFXPXW
hB7yjrv1s1AzAlmm9fhNqXnBHh8ERvNEbujdwbg3chf/kjeVAbEOCtud+ybOqBkF
xQEHoeuXgIsvyUSJh4x2zyxxwGI+yhTDfslJHDoIJBbSQSpGHULornP94l1LSmGV
nsTdk12H+cmDhQz8FVZqsDTb3icfMmTAcQb5Bkqd3bKf1D1iuaNr26UB6g3+FsZv
kx4OOg7HCCV7S2SHptQ2teH/Pmq18A3CL/pGJZdPGmEUe/xCSqGuJDqA3qKDtCje
Isn3ypBuqFpa5CzXx5DDFwI6y/fEgBvv5dDv8HgheFUG9umjRmMKuwrbtFDTTXVi
w+lDd6J1A1mCqpwYAqiSrBPQKkhfqXosxFzztGYux8RNod3jncAPDl7N8sRVz3xP
+mqKTvivYdFRJIiIlq+gnWGh5SP1BJTqVIWjCugCS1CME9AS9shbqDblVJV9oHvd
acS66wjq3KyEQQSOIYQKhuo0gm4ETtIBuTMtZKkB0o2tGvjog77ULrvEGx0IFE9/
tGjXMpkQjCci9H76loMnQwxsftyL7LbDKXR8pb+HAwdsLk8vKTuvmmSeCVEnh90h
mj/xkqbrCuaGnYrdGZHtCYP4o/PxEDuIBkHNYLWGRVFwVXBjiWY9O60ksR9GbQBY
0QORaOf9Ijiol22E2HPfNt+urMKsj7N+THVO3BG2xzLZ9M4cFU/x1qM/H4zoIlbJ
CVbFd3BijB4YnH0un8xWp8S78GEtIGF3d1pSkJK0aF4V0MTC0f6mcjzn7E1y8vAy
ML+RZEB1bIfjC6dc54L/hpZy87B+a3udxYKgXEgHeYLK3TNLkKZ8YZHp4S0vXNPM
NOBD+kuD9xCCMP/9sFTiXP1arF/j0bC2EZqgExWfyWKyUyYOQLxYaeOx/DN0r/ru
VBX3wcuh8QtoRxSkNMQvS1teiYWZEy9o+CiwWwsjt/t55vABo6FOVOGkbzCN9Q+t
hGhJPJ9sy/FquFCEZBOJu3AMVJmkMOvHzxXOWSCDAJxDA610FZNqSqI3FjDc0hKd
Wwh1HA+VeRS/7T9mkb9+pdX8P6E49PKrK5VtbNPVjQwnuYjlJqqq5bbFKqi6+ScZ
YpiPUXiUSEaHLT80sXI0uU/Ccs4H47lx2c++0pQN7oHePiNPcKvpOes2dlnrwjXt
PV7ALW6YqhIoG46GbkoEQSzGUroB7mKgQu4tbi8RmOsWnASGipybxKblvzu1IEeG
ZT5TAuFujkgQjKj1QGcUGG84nusqvOInB8pxxkyyoMzmQdTS1sNGe8yzfGQyoQrq
KMa/GXReo2m5tGRoSX9NsNZPBcJlgeIjZOEXNJV76CTfW/wSacsqRjUSTS7zaqvX
TQAD0uGVfhvgSeyvpqM06cIVnDccQaMryaLTsVqyVrtrpqXp0CHlzOtYvpDvYexG
pRyTNFeShNsXqfTJzF35sBjxHI0vHVryXPz9YhQ+lXhQQsM6pmuHC+WwANCpllsU
h84hXNh8CWBWpSZIBTnRQbqd7kSKQuxG22/jZEwjLfJczYJxaJn7xSc/ANZlSvk6
E+Kes1/xX/S3fJPFxbBSQS1WOvUsm/RbYMNqNqe/xrinti9uIV3Tsy6VcCelN4sr
6FIgrBlin0lSyadxZ707Kiz7jcqLzvlgx5l9VoiOXwl5yra9X5Lq3Aj0cjXZLvS/
RUASC8d08ni83XwWMafdtbO1lZD4WVniA69ykJo2FXPVe6cHIgtKMCpSUaAuqDJP
h2LxfE0+lkSLVCRvcZHr3OwTt+cl1ocA6F8Qa7vj3wWnlzPCRYuPDRy0+cdr/qcI
6+SpqZR4IU9SAvArA6KdRTXxGa2Ms/WjnqWSQ0lEW8a03hfoWgYJVFtQyKkhyqmh
eF99ebw5oI5BBl2pBoJNfFiL/qc/9vG5WcuJSinfpD979ycRkM1h9Ycc2s/tSO/w
5Ku859VCpzTXEJFeMttUGtm3UaT3CSE6bypbGQRMLnGs/aoAdDOnhAPS2gM0Q9T9
WF+A0RkZdNIDKpUFTsGWkL//v4cpWs2uux5/LP8L2Dro5xR2glQwHSAiahbvD4HU
TQ1GQmvo9X6+4jzX5w6o8RttCK66m0MzvUiGVqMXaYdysN1tTOX8Y0wSIkMOF/qS
f4TKIMY5vnqLsBA3sjP+9UgOlEX/XLDZIU5yeH5UZkohe+29OnOkydpBECFXcuHe
9Mafco3hU/+gl4E/INKtQ8CpuTAseS8Qrxj7ExzVQV7mN9Lv0yI0qHZejOt4Un3V
WlJhW1vq3fO5663IaNWyW2OS+jVgJs/ilwI+Hiz3MHIXhsr9C+UYdyuuDOJBGGWL
dm7zVp/3C1Y1NCWon0DSZ4844YSg9tKgjHicabMnhqLJLW49+TAbf3DHokp1hTdG
iXm4dw2eMhFaqcZCSZNCcKzuP+KSoHGNhdPSIC2Nnq0afIddqYj4+TWGjIUCo6qZ
ks5WRgbRbPYY0nCdbIxhdHDapV1lqA6c7u0ZxetCRF/Os30J1SC7Lm3oIfZp44am
pNtuTSA+z1TQ9vgZeLjohDlSb8XMSb3eoQeP9UW0L474rsvQRa3ecOyZQPR0ez1H
4wLicgxAih1VG25Mu6osoSJFXkmpyUopbJRsB6r/E/CRzKSyRkXz37WlEYrRM2TV
2uia7QLekDP4vwnBIJW8hwfXOZVvePYdSCGUE0KfRBR6GsiAq8lQx4qPPkbFmZ3o
xkTs19PaMya/WShUMYmmVJbaikUeRHuJpTL7I4xFJfTvDXqAeO7qK4yE4lIkLNd8
DGCNXsGC7B5py3ap4IshWWI872XqS0zY46DL0GwX1K8CXvyZI+iEXNScdb6kohAf
6LVbDOeQSBTdUH9PSQ1xJOK39577XrHAXLxVhErlEJaCCgFrEJ60H2qCQNgHPdBD
UQlWZuulMN6rpeY+i4NzEZTNORUGEj4v64YSfsa0aPiZvARBh0HEliX1T6NGPNPp
p2zDNhlWLd+Q1x/FnQLCaH9Ky7Oidf8ewrNGjEtlk9kjbySeo/YpXbgmQJCSBuNN
0VuaJCmbl7idPK5oZLgbf/FRFsgWgHgiiczlLuRrMkycWPM7ngMuBIxja6bDqy/7
fMmfAawdIu0MpLTYFDPSDjVZjQT2DXIyZOVn2KsDaVPuGPxU9HoGarlYoMUoG68f
ma/nM89E5SIwrSrBLuJy+N0u6TJ/wu8D1NLUEZ5DQn2DEp5LevCEJhMY0qWWXDZw
RkPG9tAprP6VbJIA+s6Ua29CGPr9lwIWDAgjSBEQKz8mw+UOzDOrbhFCYf2kEVS6
tij0/sdNZ4hvGjogymxn/xbNefPWKZIAQ8SNDpu24pQhCMPJ5zYmJ1yrXfs7d3Vx
2Q290ZxYi4R6+ajHIXD0NL5xtuVGgmWmrr27fxgqDNtrF04AYVqQmsCvCZvMFhpz
SpZo5m3+l6MKZrz2ag78E4lgv10g/msClrIqed1CSqayaGp0B6or8KiwSDksPIL4
pGesEa6QhE75eE2nY8Ac0HG2+xtH3JzWPWwnas+xT/wTFmuFCXR8civsGgVNzpP7
yZldovzFdvIyQI7zYqTZJSKthv5UXaa82V8oX3r1GZQjc10WwrAJ0865hNk9iaWC
zASaOQYP80+XKFpqqudi9UBhFFhSN99a6CiAMstsUn7Kzdci1RJyW4KEwtSsLerx
dByFqfP/XTpLPBi2gUhcE479BwleN6krslpNYbFRihwbvBDZlTk2A9UZELHHvgwz
kuT2nEvKV1F97/MW9Y55vDox2V6j0g15RJXgXlEPeP3cFocQ8nYerizxAjGQwWd6
2Ozwi525E7QcnLywssjhdPUwXXeATTb+FpwsDc2jYWE3jryJijd2LdIK3SbVe5Kh
lJnkXuUU/qKrj8uwQaUDcKMiEkW3dhTFmLwg96csaImZOlSxY+YkrdMuxEkM+Wo+
4K4IlOIUyLsXMb0X3IAiASzEBsI8dIlv8oMeTfeaeUn1ILNlUTCDduo8jQmjAEgI
onyaO5nFm+4m0pv4qZb3Fs1gHypb9KIAM8gkgREXtsUdzcy+Wxp5DUjHVgWq2k8J
adPUHDttDRQqCZptUUET+mST6n6HI510VUqM/gZ6pX0dSX0S0qTPPvGDfCFDfxXL
by061y5BrVsRCaqkGTEbnX1u49UHG60HeaEfP/jUbMbJPDhiPe4EAOK6PbnrSN7F
axx+3i4UBGirkDbyTIDfaLWhJVg9QrQbRp3m+9wZnQXh3udHVStDYKYcuAEd828M
5RxyJNGpd9z2kUbqZG/w+2TaEIUY45pu4JSCLPd2FnKmAkEGLhvxpVcVo0hY33Xh
5b9aFOL80kbHx7I1phUN2xoHce1Jf8J0o2UlD1Uc/y7q0tI5M6lOA+Ga+jmLWku8
EgTfSnIPESu2eaTKmP6HlrozC5ZJIm9k/zKwE1kmEhdNFqG4q6/A86qLGx0dJI0B
IZB1ljsCyXg0gbp9W59bpiP+Q4NABQRsGw/DkSAHICrlmelO4RaM7GwMt8hCVVXX
2SoAWJRCZL/aqaRqYsr7TKZaE9Q7aTjxkne2PAdzKbQJTagKm4TxMMX3YRCKqTfg
3LtG5sH/ucxXOT/2YZof5hfWaHRKLWwc8ldeofrDjkuOW/pcJgWfcAPTzPlb88oZ
2L4qABB2gNXJvxwn/vyiF/8NxCssiciRtxsVtkflAWHjsv00HB4JQljZrO+kcoqH
9DJBbhf/dbfd41e2sEQaQ+42knmhMH4N3PfCLoGicYGY/9wbmLNQUZsUk2A11a++
+nBdFxIOcP04oIOutCtT0sqtSYOp8LRcXlmqJwFK8E4a+JJl40uQbymXZD3v3MmT
g+5pUygClYV1VXm0RYg7u43MRyr5+hdKEWd9ehdHLaL4iTIW5p1Vm0bDrXJAtxMz
cOAN4QCruC6GORrxKgNFh10OvFIS+OZCFdMs8hNPezB987Su7V67OR98t/QaidJ3
spPR7vUgE58T7gB0C093nDdDGFSORgRMK2Fa1TSrX4r/dbKVUW/0CCKTQZDLh50q
cCva5hJHE4E6fAmDWOia+7DnUdDDvYQ3XmTw9qp8VGtwGsb1qzebHDWMONbIxcBn
1PupNgEpnj+2IAPK/CFBzaZS+7ukMgGN5YPpSmfxSPV0kRMCCIe+Wx5yeK8OjLRF
qdkmtOzFDXMYSVaqFOFw9cHQBjP0sPyiVo2ResYPGir6ML5U6LqWYnJdKJjPG4MZ
Fe2ODyqNw5vZoT66wbPCmVQKg+dvKQqAEKDyqN8j1uqhOhPKVehdQa/n2sLWVr6L
MmmM/AGf3MZkOkn/T9m47QjWRTz2o8C7ualzhkc7Z4zfUVAgCK1XDWWMOqwhEqqs
ZQaMCnLjFsugGvNEOo++2vtyjmygP0sfz6K9FYt8IikoQTf+ttO86nYJ764ZqlMC
nz/uz9+lVvjK85lZoinQP9U2Dbz6m+603GyFGd1t8gKI7TFzIAEetcZYxP2hnOns
iczqdou8Dm1DV9q3PrBJBGbjwBj8cNcm9ri8KRozuzRRJIcfGokXUbChlcafH9A4
7zalbwDaEg562l4/Hfg1whB0WlDyPQ9Ft5WlK5bx+XsKsXDgBE98O9Mj5TMIlfEw
ivs08wGQG5h10sc2BinpbI1wwtu5pkBly0ecZcdSotLKopqDRP5gdbtEe9sdGq/p
C0UOC7JsPDeN5jEGf6psWR15/XhZHDW9V8ntZCUmnEUb4B7Na7snUcbRVuEfwIRg
TpJuOfQ4ayOTYhQS6Vq4kX+wOyexvdRrnL2Rbh1zhj0h69gcXTD+9vyHaCjJjc3w
S5L5V3MoU7tIU4yHnggyJU4LLVMlGj9enGzbwoximjDvwgOu29M/QnUNz95QZxKi
g2KUGy+ST1tFfLEkogyR+1omqNaRfUBR8ymQHBtOyd8iTuMSSikzEaa5a9YjTbX+
Kx1atIsMrPd8gDyzEnc8BZB3vxGRtLgUR2x6svYkKOTv7Sb96ppNYFTAXXwt9Nt6
Z/0mUNpecx3IR4rbmpX3WmotTmzCS+kYpYkDtrybdjTYA3Xo43RqcN/ZLpRrDZQ6
aVBnVoAuxuPu840L7kQQez0vR4hBwzvU8eSeYaj305Slrmyf4RxA83bClKXnFh2p
igekkT0BC9PF8UBwCVSQJIL+LEpJvscUuQEEprV9bmmY84dDcTI0MtSbmnUBAVE2
yahHw/719kNeTPl/djcfhl9BhgzAPXFkQPFtTNsNFi1YVLeGMDbmFSToOOIF0mv5
acuocKkO1/g51GKjGaZ2oagIjI0o/jNjexK/qzLpqRokGc++nRF+ahp5VGGVzqDl
O5eppfD97BOLkrVXnoQp1Utv/aG0HZrIBVbANJCqlKh+1aeiDFV7/bOukTAq+DeJ
mS+oS78iq0EHnFvKI+TYEQhXDSIHAw6Mkus6eNkTD4/2XvhoFy33j5iZG06WOmKl
ab7G6MscFnw0zhtbTnPn4r4j/cy2nw1dBbS+5TJxUfdhwzopSc5pQgecaCCT91/r
FR2hj7voStykY6eR9x1jSgSONWin0TCR0yLwOo8jzS48Xpa9spRT2CjgTcrDL3DZ
sJ7gjFaKYzJkWS9bNGmJpJMBvTqrmwDpM2SxXVev9WLgNnyI0Z7rBGwpbQ57sI9s
4VjZzpXmfd1WAa5EpqXlsfVuQgYt3qfBG6LRBZqyo7+J6ZHhWxtd9MPZF/28+Fnm
PT8rvJzl3L62iMjFPQlfQDiwkztsxpl2ZPK9mVn/fzl8y5bb/8Nvkk7a9dyGC6p2
D7Xc9IkKwjlQ0SKoig4X7adF9tSTy3Roq41GauhKA9YP5drfLycWRj9G+fMmI1iK
2Yz2kp65bIF+DXrWNqk2iWtq+XOk0rQ4v8uxrO5M3oSDW1WGL3vBaSPDikBb2s3x
XQUKd/SEcdsehjFf2nmRcqdd/qYiWQxJqncPcfOt2nvEh+l+O94b3YFp/xyqtnOX
fGSE5hewjK4pMOKNSWs+RBDtXaTK/J+HOVKiivgmD4U/R7TPQFACeEIwP7KEuq7A
bWjOf2ZtqSZKQBk8mD4u6UN+IDf635Qxv3YEH+akH3cC56OwRFMej9Pn9eAkHcwL
rwjhb2YT38rh4fj6jLB27zimc+9HPc7PNkXbsKAdX7LKOuE010D2xVQp8XUxNT0v
v2MQgWrsEtPKzjHFtQwgVz6co06Nd+m4wjeqBKUdOwH1Z3swLYc5pl0NQh4Avh3j
65Vg1sEJ1TK6KMUg4OhGfukw6FQOHKtYkcHNTMFkeV449+jPoq5kwRrj9qE83I6/
d1wUS4wwEhZ57wCAG7iP9S+zAadDHVtTdvUBmQTNyoFhwZYzzuKEh3QqJuqB3heP
uOCz21GHlTsusDLqeX7f1LCoKCpxZuypYEEaiPQwqJE4Xx6UH4EzdIbhtnMJZxEi
p33pLEQT5R9PRE8yhJrW4A==
`pragma protect end_protected
endmodule
