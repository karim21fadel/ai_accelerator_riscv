// Copyright 2017 ETH Zurich and University of Bologna.
// Copyright and related rights are licensed under the Solderpad Hardware
// License, Version 0.51 (the “License”); you may not use this file except in
// compliance with the License.  You may obtain a copy of the License at
// http://solderpad.org/licenses/SHL-0.51. Unless required by applicable law
// or agreed to in writing, software, hardware and materials distributed under
// this License is distributed on an “AS IS” BASIS, WITHOUT WARRANTIES OR
// CONDITIONS OF ANY KIND, either express or implied. See the License for the
// specific language governing permissions and limitations under the License.

module boot_code
(
    input  logic        CLK,
    input  logic        RSTN,

    input  logic        CSN,
    input  logic [9:0]  A,
    output logic [31:0] Q
  );

  const logic [31:0] mem[548] = {
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h0100006F,
    32'h0100006F,
    32'h0080006F,
    32'h0040006F,
    32'h0000006F,
    32'h00000093,
    32'h00008113,
    32'h00008193,
    32'h00008213,
    32'h00008293,
    32'h00008313,
    32'h00008393,
    32'h00008413,
    32'h00008493,
    32'h00008513,
    32'h00008593,
    32'h00008613,
    32'h00008693,
    32'h00008713,
    32'h00008793,
    32'h00008813,
    32'h00008893,
    32'h00008913,
    32'h00008993,
    32'h00008A13,
    32'h00008A93,
    32'h00008B13,
    32'h00008B93,
    32'h00008C13,
    32'h00008C93,
    32'h00008D13,
    32'h00008D93,
    32'h00008E13,
    32'h00008E93,
    32'h00008F13,
    32'h00008F93,
    32'h00100117,
    32'hEF410113,
    32'h00000D17,
    32'h234D0D13,
    32'h00000D97,
    32'h22CD8D93,
    32'h01BD5863,
    32'h000D2023,
    32'h004D0D13,
    32'hFFADDCE3,
    32'h00000513,
    32'h00000593,
    32'h014000EF,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h45051141,
    32'h00EFC606,
    32'h45850420,
    32'h00EF4501,
    32'h67850D60,
    32'hBB878793,
    32'h0037C0FB,
    32'h00010001,
    32'h27B74711,
    32'hC3D81A10,
    32'h1A1077B7,
    32'h0007A423,
    32'h08000793,
    32'h00078067,
    32'h00010001,
    32'h20830001,
    32'h450100C1,
    32'h80820141,
    32'hFF010113,
    32'h00812423,
    32'h00000593,
    32'h00050413,
    32'h00F00513,
    32'h00112623,
    32'h0E0000EF,
    32'h00000593,
    32'h00E00513,
    32'h0D4000EF,
    32'h00000593,
    32'h00D00513,
    32'h0C8000EF,
    32'h00000593,
    32'h00C00513,
    32'h0BC000EF,
    32'h04805663,
    32'h00000593,
    32'h01000513,
    32'h0AC000EF,
    32'h02142E63,
    32'h00000593,
    32'h00B00513,
    32'h09C000EF,
    32'h02242663,
    32'h00000593,
    32'h00000513,
    32'h08C000EF,
    32'h00342E63,
    32'h00C12083,
    32'h00812403,
    32'h00000593,
    32'h00100513,
    32'h01010113,
    32'h0700006F,
    32'h00C12083,
    32'h00812403,
    32'h01010113,
    32'h00008067,
    32'h1A107737,
    32'h00470713,
    32'h00072603,
    32'h1A1007B7,
    32'hC0164633,
    32'h00C72023,
    32'h00478693,
    32'h00C78513,
    32'h0085D813,
    32'h08300713,
    32'h0FF5F593,
    32'h00E52023,
    32'h0106A023,
    32'h0A700713,
    32'h00B7A42B,
    32'h00E7A023,
    32'h00300793,
    32'h00F52023,
    32'h0006A783,
    32'h0F07F793,
    32'hC017C7B3,
    32'h00F6A023,
    32'h00008067,
    32'h1A1076B7,
    32'h0006A783,
    32'hFF010113,
    32'h00F12623,
    32'h00100793,
    32'h00A797B3,
    32'h00C12703,
    32'hFFF7C793,
    32'h00E7F7B3,
    32'h00F12623,
    32'h00C12783,
    32'h00A595B3,
    32'h00F5E533,
    32'h00A12623,
    32'h00C12783,
    32'h00F6A023,
    32'h01010113,
    32'h00008067,
    32'h00000010,
    32'h00000000,
    32'h00527A01,
    32'h01010401,
    32'h00020D1B,
    32'h00000014,
    32'h00000018,
    32'hFFFFFE5C,
    32'h00000048,
    32'h100E4200,
    32'h7F011144,
    32'h00000018,
    32'h00000030,
    32'hFFFFFE8C,
    32'h0000009C,
    32'h100E4400,
    32'h7E081148,
    32'h7F01114C,
    32'h00000010,
    32'h0000004C,
    32'hFFFFFF0C,
    32'h0000005C,
    32'h00000000,
    32'h00000010,
    32'h00000060,
    32'hFFFFFF54,
    32'h00000048,
    32'h100E4C00,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000};

  logic [9:0] A_Q;

  always_ff @(posedge CLK, negedge RSTN)
  begin
    if (~RSTN)
      A_Q <= '0;
    else
      if (~CSN)
        A_Q <= A;
  end

  assign Q = mem[A_Q];

endmodule