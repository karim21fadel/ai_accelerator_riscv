`pragma protect begin_protected
`pragma protect author = "MED"
`pragma protect author_info = "VirtuaLAB"
`pragma protect encrypt_agent = "RTLC VELOCE", encrypt_agent_info = "1.5"
`pragma protect key_keyowner = "Mentor Graphics Corporation"
`pragma protect key_keyname =  "MGC-VERIF-SIM-RSA-1"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype =  "base64")
`pragma protect key_block
PL7ByG5e93DSTzOTouBv8/8XbksTYZ30QNyHZ+RDB6x2oiR+VnIw+yDan4ZTul9V
wiCZhbaCYa6JmBJvEp8YRfY9mJxHdyIQl125V1QIMwckTnLeUZHSjGw7ILmG0JmT
7dH1mSS5SPtRIYKLZrFfVNeUTDulihR+dls+9e8HLqA=
`pragma protect key_keyowner = "Mentor Graphics Corporation"
`pragma protect key_keyname =  "MGC-VELOCE-RSA"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype =  "base64")
`pragma protect key_block
tkdTIFnU1K2Tqsc9uzRgxIsIgjlxIpzX5jdQvpV+xRd8yHcLS7yirfi89g3bQJ8Q
5DBGAkN6C5hJ9OaSaQEtBYfHQ1hNoh3ncLSTGzOddYNbWzotFWwqeJfva3LOqK5X
3hl97KWoVVAVqzC2mwlbkdII/M8kC8eltJt3AfUcM8E=
`pragma protect data_method =  "aes128-cbc"
`pragma protect encoding = ( enctype =  "base64" )
`pragma protect data_block
XMfHdmFmTqCWCArz8t/U6yfAiJScEAjuGqu4PUJ63IiAjVfMXfG80FZYvube4Epu
niwcLmCXTHJpSJZ6lKzfvDnN5C90g/llvTA7PfM7Wulij5+xCmfFTiV9vD+R5OKx
E/Whmjb88bMgJWjQrFEnZ8fTnXOA/bD0DQl34Iku5uokmA7N+r5ui123tEhPtdYG
KtUUWyV91ryRGLbm4L9EyqHhY12H4zs9mCjbXtXweAAjg0Njn8KfsIPBRGu6YFmp
Dt0z7Gf1FEbX+EgmZBnOj3pMjSmcIsE8m3P9PNRIGPpR+mLlrYMqSykWSfvUejw1
ysSkrRo+Wh1EpDaABtD/CmpIII0UPKGJvM/J3DtiNAr7doqdnctbMCZ1Jf37vQeP
lypIoQzGMgortbADgx+8uHNn5qulHSeMB3YK/9mBmTS6G06lbjBW3akU4AWUN5aL
cMoYzk7ID7kLH7ajClnfDVsULP4sQF12UNiTQ3GwimOJ7FpQwAr8c98agUhlHUKg
iUx7D1E7Gqy32Rodql+bTgndEjzmu/mbjYyfrEdS8yNCrhhGqIjV/1Tkm8rr5i0f
TbzoqBQG9fqBLFuu/RUCPGzyBtVjN0mOiw++anyDRYI40kFigqlzXsIEgfGrXWAT
2DSow/rYL9HvTrR9YqyOBMed3qt9rq3ck4SMvk8CqftmO/XO5dn8grXxMCmWLg0j
lS8sVaHVkcyM8AycdTpD9XvpSF4twO8BfzyKbz/nQy5p+SpcDiYggEbX2Oz9qThs
IB6FjkwgLIEaNI/aoj83zWpAR7/eLUEuFPnrI60RYIt5XeCdrfmRJ0xozyZOqNSp
iIEX1SIvOTPyARTRwM0EawbfyPYUsRmbvIQ7iGyp2GPfL4SWJKYrH3AHz2giQTNg
MibxH8IOAJv2rT1Yb9XYwNHAjCi8Vdo6A5/PXydwl7IIu483QaQESI+/h39tVjy8
t6FWFtx7bCKF8tIqy6AsPCJJaLWUU8TpAQJ3euRGlFXkZ96ckveu6gwJomputYoL
ZVo5uSRxu6/rfxJYiKu8lLvUgpNvhvvzCU3Yn9B/qMEEExNeFR8bmMbB/0bRuXXo
3cDuMy2CYjTEoiHOmKXkLJeJarFmrbcsAay4cctuJPKRAclG0tuz2kMXAue0Zas4
YBYhwq03qDbs7oNn2spYU1HHGn1I/Szlc6XqEsjJ+Cnq1ENCDhS/O11MHRwtpKtB
mKX9RT5FFV12kz5vgzNHcKzX1o+8ziXwmRh9xrIGCSCQC0vcnS+NIcTdUXkld+NQ
HhGFuIagg5Gz333q11AihPlDjFZ/Wnwp8Ed5TbnWRsw8gB5h3sq/k12F+vHEL+Uj
7P5lcqfWK+tupy6hnyw8fqnUa/vIroM5M4sh8uIT0igURxuCa04gpCTAGfkS13YQ
XULZFmer0PinLtUTOkJagxQpPc44UEKYxk1pmIR7hOEviHk/LjcwIRfqRjBN5OIt
qKpcaDRNUVN+fEgldcdoESFDf6QGf4Ah2VYLvyiNfTGQMl+ZSV2+Y6UGemlbBxDa
qZmOVef986/kRsRqwIeR8MNLqm1C16EVztEmewy1ju6XQqpBftVRz3gor46U/Qza
Ml0hrPypRGx1KVXkqvHiSy/Sq8yhLxLpl1X5opq1Sv8IYdRCuUfaMLkO+rw5xWFq
Ek7pxjVeQ+KgZrQn3FIsmvofmVND79HcGvdarz3WKpjrOPUJP7iIaNAlo2KoSHLg
3RoMH0+opKncdZKiq72U304vg2KCmXvUBTNFT/jJdVI1EpfSaYBmoj9V0oBxbcYL
usGXdjrOA7KTNAsit72T0H45IUXKOam16JyWgDOy4Z5s6vLbAqTfW1YlJWh+Roi0
ylllnz91Q9RyELfHewSGvpT3/kJQIB8LO747iX4lWsBJWJLLTMKLnTdXobkxNuSP
ac6fzWuevwUfDzSIPq4WqNwLRJCOZNvofC9ziFDwyClvpQrFOwOv31CAzUDoTWS4
hFgsDm00FoDR3U8dfCzC/FHrBf85UQ6HR1O3/SLF1Vxs8fWvQm7nfmMHBb325ZY7
27y16KWisUmeBtRpjfjSImcvGKUzYHHEqFgn9uGDNZB1guvTwop991lVm2UXBKCy
Orzm8qESZeyUFf/qHdH8/NYZzEt4Hxej3vDcrQ4RjXvTvUzdcMgC9izHNphIN2In
0XPrxDwpFvGz05z19le/WUghdc7roatWrmr68bHxtGbFl5dvknT9qcRZezfswDOv
KmYSMBPCW4ewz3o9mt5IJHn5wi2pejC1Ay1RGTG+RwO0Ty70h1el8q+ocvKocUQZ
lDK3ozpE56nIUPfxIOpAP3yH28+/4RCux8EkFB01G72kirxwTQAerniywTkSDYyN
aiyo5rNXodM5xEjkYYIvl2Q+OEqfsjCSDqKNfmG6VWGiJkA1tQhrjfa8p4e1HHU9
ROtp87OEaqpaJ3/VYVDeMOluomNSVYO5ctwBE7D1tWcFVWWDHx8dMqpXFPIw04jH
NCQ22OB4ClQxDa2BDa9fOwQ10Z6WZa18/CDEBOg5riluI89BhlVEcKmcqWIaVh5C
azciBHSXzf6WXy/S1bwuZkHFDj2cG1G8HAM81D9mb674hG/z7jIjWK/xeAzGb3d+
DnQcW9ZFZrYcDJMb8ptZ8Mb4rbIoMUgKeTjh3VSifhlnS4tf4PSGq7aa3PKN8UDe
46/DMH/tx2ww23EALFbW/ql7PrJkLLY+BGIxpsaYKHo3BhCdJkAWAREx8UJWvb6N
mu6DI7fxr+tO6RiNpIlHoasJORQ8r8UreaixMGD6FzTvcFIzVQ56Vp40/32d1SCx
0+RSPoDYD2P+QrGhBhcyjVp3WCj8L4UYDBn/223lEOPOpLT+Sg9B1B6XyOsCilPl
je1Bv4JQ+dDnh3fmtMEYUMITLpaHnjG2Vp3oD15AfqVsMJjTQ1qDsMN77qG+Fv8Y
IUmCRItUcXvmm9w8BpeqzNCTspYXNC4yrER85zqgNGgkI9DemyRGa2njdlUB8sNW
EyHDTODsftbjxmqSntAnIS7aaukNWA1ZwkSD/tv5vfuSaYUuXfd65jmQ6wjhRkbX
4FIGPxB4ErYCKOt0bM+nl1n+VhWYxvQ3Y1+7T19LUhv4K4onEjXCXbUGJPKPcq9d
kQBIZg6sDJQ++isbQruvOptbuoeXaa5RxYrSoU+KmCMmoqGJpcZO61/RENibn2gc
RXXv7rjoErsklzih1mEnF3jmiOt1RN84Cd1466zIiJ/I1LumGwBK0zTiHZr6UFrN
/2+p0rL6JD9IRiQm1X8cEnjClfUSr4yeMYwKPq77Gkzr1gLpxly9kQykyNk++xuC
R/6DJ4w46M4bQvaN1ASp/ZLsWiPG7xYJJ8dG54/Eq1Wugf7HSmX4L93kc9R0n5VA
LAO5/HTiLFUo7/5/EgKmNmWYs/8Sc9kYkshKMD/w/eNpYamte2M3B1JkaNmK4RQm
UVOqINjgjqghpRVmdGH/uKQFwN5bU7LNr4EWiVnaYzkNhTtzf4VaweccPit8aSqB
EpeVsfFJWe24mgkyKkQXwd/b/u4/adTu0Ds0hTrCeAK6c1o43vaZBFEVctmIKl3v
EnShPzVFpgaLgAeiI37zNffRsMFLSmiUYtW/DKF9ObtxivR30hMaYD0lNi8Rz2NO
8n+ccQ98/4TdlARQjJDkNgLZGwiSY4sDh1xVFnrHlDF0c5bLcsbVs5ei4JqtaPM9
3MiRCKnWm+qrmdfjNWPtb/iANgsPrizU3vx5wb9apHcX+ETY8DzvTWC1bkPlBCXQ
L968BUmqcQLYZkxsD4TBOAZMUffO2YeuzFL7QxH3dOkIpDHonyy484kkvNDCl0M1
NnF3UmkXKolYljAQPWghubmQfZd6o7JCFeZo9LNTI8qxb/DWbNljtB3hY7xbFdio
7Nhl4a0dFKDIyzvE6f3XSWBbgGc7ezkaaSIStukurQlA6XExbcN3/abfiB1VRhtC
h3UUsegdaa1muHjzqJEQq6zTIR/BCfKAZkvt+nXbQVK12AhL9lXvHYsCJ5p9xi/N
3qmzNlmVm1Ux1QVNX2Enc+VNrU3FKOyqaNsK4bxqBQwjmoWhbgWJOCqzYjyNCB7r
AB5SXMvOeYzXVhpMV5tbyPkyU7VVe0PQr/3gz/yZ74aAQxLzPKJCqWVntF/naNxL
DXSzJgqnixdBxORuLTvMaS/oJNVPyF0454ZSZUq0GGG2Gf7AIKtVvEaBvg5g0wG1
ZjLO3qP1FijOQLZbYcus8yXzg7JpVf7PCgi4VTLPHwavWy7rhQ43Eu4ewdGdftdh
2I+NTdG2YQC4VEhIdWPIRQkzNuZcJhYezw5xqoV5uBkGFOGC1JeXC67YlbdPVoSm
1jGusDRjT7+lfst2HH4xImOdyoB4wcgcUiRpMOdb9HoWgiNGP+5mswnfqRQYeXT7
91RgXatG/HeYaO2jFO3K+89ssdP3UGIWl9/7XuZ2Ger46m2hvV6l2CNlu7eW0ZJ0
TI6KOtQys9cSwQR1kFJrwSb9u7bTJYkdtKSaHKCoFcS7tRrq/MA4Xm5p9NRD8xpl
aqZ69MjHWxDNAqtzb/k+tyOiTPwqM9cI2Y1py3rGxr1F2yGcX7KVHD1s0HtL3an3
x4AHWfK7ghpKpiZEeSGSX1RzTCrgfgnA4YWd49d4s82hOA32VMXO9pq5Y+/hvsYI
aslQ/0FEhzxO+Gk1Cb9T8PH1iHkjvk18ZvFvhSciwzf/8/c15ifPavEXecz7f/WU
kvixG8XN/CSiPNuZibl8mMHshF0QvWuJ7hUXg/z0IQqFZYfVfw6BydFJEy24aDe/
E8LY4ddNX2Y0e0YWYXmiCMf0/35Dh60LTTXQKvg1qSW1COobEzL3mG6Cmy2hoQcc
J5Rr9+qT+AGC2PbSnQUdM0/cxSmJUTbSLRJSJi1HWCUR2YGi4gUYtNvqZ004+LcI
uGEdYe2uXLTOoWpZP8DPJQNKdHZRIhVaPe3hezkqO6I2tBGPAHFumq+Hmd3Tn+52
PlZ/Z1V0GFxzFlOPb14thO9AApe4A5OrlsX4z3wApIAFDX/t4A7m4o8LPQ99TdMP
S4al4Ak6rzqrp0NQMOsjwuJJb85taYmS2jcHPWWxbEayrRtligZT7TZeS4OE2bgL
AT947cMNUY9WBGO6jYrGrL13wnCCMIAZHKgEoJXkNHGdOEj99vOAZl09YqFaoTRv
Bq4+XGKPtDMkvhJZa+kQHr5zORlX00o4wrwBfu1/tJlRKI7rbjZ9Bx9wcvahOurO
/x2HGc7YRXYdJ86UuFYtQgLuAB87K3z2oazhIOC+5I1WaH4nymzyD+gq3jiX24LP
iTqj6YCtvr88eruHN0L70z8ijsMr1p+3QilnmDMIj9SK6BtSE9mWvwuSZ1ZpffyK
to/f1qAyK0UpVYIMGtBqN8Sl41vxMuo8wnex0iycK+cp/nnpq7gvMmPuGXW8/1ki
0jbYUlhM9zN51B6Rw092w76rn0Yn2VS7EP3D+3ort75YLA37IeAyH7kr2axSP0dL
YLgVPPLzPBM+L3QyUD2/VkCKLzykrSAHv2gLx/6z3OF8btK8oWQ8WO0JZv3sHopl
K0mj6ADcQDckIudO92SRXAY9o1YoZm6ksohRozaM/3wOYDgpQ3yWTj0JX7yK8OPw
Pl+RogtL/zn6kzanL1Rx9+HwefAhm4pGEZr9iRXDUj/GSDJ644S24esHhjv4+bVb
yTgnKOQb6jjdHJbK42GHPq150EOryFU1FrDcH+h94EyxnPmHjM2a0+1O028uyC/T
DEsjgFL4aHlnxe+X3iqqr2+mYfPZ074gZQc2Bo/mtmh37eNGbmkTfTyEEAbH1AGC
0kgWP95tHw61Hmv2uWslmdHyUDZMm38BE41k824+CzMYmhCMg5N1sC7QolfBCPST
+7FQzqNIQs7/WaYxnY45R4VbsQVp5ADVRYat80HZLaG268zvZXnm6M/eOYiKLAmv
jL8JSYTAdQT9lghjqk71eh2LPR10w3V6nI9vU7CfJzb/bBKbquWTEZvjcqoz/e1I
bMqPn33N3KId2QGGhYpJHq7NG/QBLZQa53bT+IgcYKJnphnun0gz1nKTUFALVG8X
YyvUHjltUlk2ToLV9+ecBrg8jTqAvHzxtnu52b61QD50F780r+bzUnAmoIP2dm6+
6+BQv1HtMCx6PefSGL1rkBRXYCyi5cEOPc7inxF+Xp5TVL7zc8dbndsf3+1/wHJX
mB94sYc/VZkFdQVAVtqhhOjEU6RqXGMJEK8quI+VNnYvAyyp3O8uYbPcXs6pQX+i
zTyDGAZy5T33jof6VFxuSxWHQbG+B449OA0v60vcsEy6v34gl+P6B1BUZwzvRe+t
JF2ARUC+tgw4VxR7OmRqSTD/tU8VpvapPsY8SXx5q+t2xGi7wRJCe+ITd7MQ5UT0
xN4WSVPhgrnPCqw3q3/x1hUVyN5LoHO2AIME7YHxiqpfdz9ViV9DXER/VGMFsmtv
zGsYf1bjt4B0+aosbcwWEyLInMJgoBiOIqt+nAK9YYKvayRGsVQh+QkU80bk/M65
zhdOXJDntL5ZNQp08U9otU3F1l+5iqMosE0OPoFvWfGLYq3SUVzXZYVfW1vX9Z90
Zk/bDl4gjTymds1w94LDmnj28W3NUho1fUglzDCIwUPYQz66PMABddqVO54aeRsg
Nn3bmuCOIbT3qleJ6B5rJKuZTd5KQg8mUkbBMWCRo7QxSvDaOLmbcKMUjxbL+Fx7
H7NCfUPSh7GXAbkFTMYncbPlUvkhtTQgFaM2n7cxgv+wsRxBQrZ83j4HM4aaeRog
FX0XiT/TaBOo1oyew1YoTkhIcSgEyH8KGCA7Xp9OFQKXEQwZL5nfnVe7hScmYhLm
hnne2oCYcUJVIv6Z/aJL36eN9wFmEHz92KHOlgGJU9360YeA+wXAoSEEQp+wDjuV
cYql2Ao8nu6OEtHoC8exjWkx47DLdJzpUZ7Le6mcmsoozUFxZYmFfj8fioqrujRj
bZDPlvr8SxX+FE0Lkk9C1mS11k9xCY4AnWceYvWEUMQtlZgM4K0wyCpEpICtMpio
tgThB+9HOXdwCVIal802v+ME0Fu0ZTSoRPMDDh48h0Iz+Luou8K/Cj+AlEz0aR/4
QuAkaHL7XhKiuD+Rv9Q+N9hask0ZMpFjKP41z9pCA6k/0vT65i+RbdAE6jhYZsUQ
vwciBJIps1/OVhqg2fijmVnkaqx062QDuUunoREt3bgfNWDY55PAbS1ls70a4WlC
wYf/VEZpzfxPIRAO6uZC499gNqfzQEPi8RkxcmDpeZ4buIk8Bkx7NlvzHEyoO0gc
tnHoKx1w5wAbMZgBCke6+T2vhHniLGhT6tsRj1EnJ5Iq222XMMNCJcQjX1xXwCKd
T2z4zKgIDDxCtpW2ppmup7qdXZzhB6UFPHbgvKJLTl2nVbboRH/SfZClJEigL6fd
dYpK+JP4BGDAWH7mlHfVHkS7EN/kf7yn76P2ybP69UUQG0IbQ39FBL6zy720QDE2
nVGkW5FoWylg2uoMCGMTb7UTHfKQl0WQGMDRZ8LoOpT3e040/6i3R2alMZFDZzJL
D3twX0qVo4ZEJk+UJv3P/jx4PXO1C7tmCxTqC2c9qJX5Kx8SsYuYB38DnBFHLzRS
2GFbx/J8GN0x7m2dktTOva/DS/62lauDwg98CQi2gz7DOYynoym8nlzHLag20vob
hsoS6ITV+60pWHOs0i1eTNNndx2vyhCbBCErm1B0fch6Lm6rlpahexCwXbx8B4ek
+aPxJ7tkCVZRsPNV0wsu45YRbjjydtSU7G3CZo7eoOLcSMMQ3cJWmHgNwwDDx9Go
iSiLTJDQZVjCfJo7k57RN4nOk7KEXPIVyhKwHPh8UCP9yoD9cRvu7qs9mPtJ7vZL
EjMQdKgkpr6sANLSJ1bTVokL6eEvH1JrZ/rkP26SRbSYicAp5hJYv2igjj+3aOg+
fUBpkQOHmYZmDSOlwScXoIjtIbRz57Y+NCflZimItWH4a0HAf+gXu26LadUGpPlh
Trpd0/bqaAbP9rPJ84gvHefBLwnT6mTX99Y+aWB88QUdBKy+xegoiaN+1CqJPEfN
bXK+ydhL2BEKbTWpTxY2YvR1XhPL7RUbQOMKV0hnyDy2XjrU4FajvyPbe+oaRFC/
RmMaT3OZiwAy3W22hRg+ta60ADFafig2l6ag4BRKw02CAl0UfnNpWa2m5z1Wwq0T
bBi0XVbJE+wrH8ORB5XX9G9eXfxwGZ8sp5YFz7owrqClb31+mgbZP52ocwZsvNcO
cbE8r24IgyTDUa74S3WVq5bKPUlPCT5g78heUXdrzvLMEyWC5Qpnb66+9x6Xdzns
cTTg+IBxiYxU2w6i0ofP7LDMMEo/EmXxp1MgeWWWBWAbctKqKDC9rkDbhdEXfMNz
QChl0wyWsKVtt5Qh/jqtkyjzfn7wIAFOgiovIDhS/hidJ4FzW2MWyM+0uUH8Ja8h
BPFzr54X6rT+6MKkYVlT2wId46Kyb28BdjGpsdpZ/wCHyH4etnNh5+jtP/c8+TNF
4zVHizl1GOsWXUb4Rh8SDZqw6t1oumtU3FTDLpoBGvSJ5PDFo0i/Cu+Ut44MNxqI
ilZMaGvruddSf8Y08PSATn+eNFldDKn4itIcLd1CDXUvyhS0+TjBzMuUWBM41Szt
WX1gZ4O/u9NoS+U9M36y4omKjETy75hptqZ/MX9qLvumI3vLnS98Es9mdcOrTixX
gJH1h9styqVH90DJHKvS+AS4DftNwQ5uF6b1Qoa7Z7iIaZwJTCZnA22FP05r+TQ7
N7v6wpCqzFUmGBu+e0SuXyq21baxzuqo2Ig/6PEAaYeu8j2BBSpCdEDP8JQeRrG5
R2SkK6wIWLoPEfItnE8sFLsrYre9Re2pS6NL3xSWPPxP5p3NUAqJ+7d0jx8Xluhm
dIoqjpQgjKbAqZl1VuVdb/33q1lDIz96obRTp2Yrs63Xk5Jf/yYVvJgdHZyZQmUO
LQi9r/SfIeTf9Tg3FgzPBhbIj7dY2fAm7KLCmTQo9vpTV49PfNe6SzrwiliadlbU
KnN7JRTgGQkfxBzc6YwIN70QZaArTj4fSrk+r43WNoqBXpyxCt6EbTv8gcdBXmAB
dpoCSf4YZSpUuNPN1RdFqLHrUSQmOPvgAm6XEKFAAlQ0CnbUtFAIyB/SlIBZYa3v
G5hWV3x9qm5SBItqrU8WvxTex5cbHYNoEXfKAuoQlcDnkjKJk+o/eK8XFdPAHC3L
ILP/18p8QIwNRFDUB/77ttOG1zxrodRFTHOnZM+M8ozH0QC1ArqCLkwPvsiezUrf
ZbUBX05kkzb2Zeyv1RklDAjf5t8x4+kLjE+BedxNmUiFj8jG5voT79GPWbb/Kz6d
C0tLNAh8DWzS8dYjyYC4zA8nW4O3p9hZeSLMbJZ0RLbeNeLJbL30Dk3G+lnLgsw/
bxBhbtoxsN4A6OHvITMdUZk/lOoXc86+t9ZV2aJUW9r7/geZA1zRJ1yo0Z6yJLy/
NA66qosBlsXT6tDi8QMul4gccngstRXwoAklXl21oVwNWNDT256FaCkn2hXcRgZO
NyolcQyPjzmCiYR3YC5ziGG3yQWD/h9w8IY9DgkGqMuMlBeLn588jp/AKd1bfZa9
Tz6Mp7oIjuEaLEgHD4Qd4wljri4sic851m4EfggYto5o3lBG9PjQDqB+Wm7UayQy
0cCkN75/sBWcCzzjKDDxrXm9ipMrR07jJoox/yFeTidI0qm1l9B+KFa5ZSHeFDJX
aEog5eMDZh3BGHWjTEfVwE+Dh8jikkfTYys52ctGFDVhXlcCxllVmBeAXzP/X5gE
J7jOAV/If39KBG1TzRTcwz91Lzh9iOQLSKjy9TnzQUMJcV6Xj2M3kkPk71O0O2hR
jmrNgpR3bpu00dlnlwihbXFZDVMZ5EINGxeupngn7o1f4csZJY6stiWBnMSXECTL
bCoM3ef7lm9m3fVw3PMH4UThqGAfvWDqMdR9Q8D2sxyb8WCNIhRYoz5J3siv3FBB
irFp08yzzw8rrcI2rcRtQIUGSr7q+4f53Qz0QEB6N8f0OX4Z4Na2vgk0Iee1uRAc
hpn7h7CZQRee/8GVaLpH6hTNQNZDSu5uxoVFjTqyAhEmcaYUoJ2xvmD5TiyUJglD
z2pMX6FvPtUKC3mnlhSMVYclQtgq441SXUF4nPu7wRJPpPAeeXjHTa5lkAxZtfd9
XXJvVOn0cGjKZNRe0E1LtA9x28KT4Tu6Ft2Ucr+jDn/neJ14JrPsAxqpuMMmH6pw
bQ1VSxjf54HeDNFS6aKkyQtXeTcq/WYPKKbx8OScOMBaSp3zlG4j4gPLMcj1r9sz
NPzrFOZDt63Jz7fzC5uN0FC+9NrPCBbkw2nvKqYJiA/OEtGAz8f8fRo7n9dWN1SH
QfEIbskmMnu3Sz00uGmRUyuSNCSCNh5HXH9zjlzgrIQJ84tdOQu3sjB0DFG2+caZ
315GVrdZEQpjj0T81yPvNHAyez1zxq+wMPzq4X5FY+NGH22pgn2bfEtBhs26kwr4
RF6dV7vDg12htIh/s24Em4DJkMqLfkCWaY5abgOT0zjg9HO6x/TU5X1jUN4vsJvB
a47ZNncyMRS8Yt7SK7Vr4R1arSUlYLJRYtDiGaMcNYU0IHUdBos4iiLilgelDmn2
z3jTDqSROFRBo5Py70cDDJoOAPq4atTVLIpySsnU4j/1mINSv9jo42WkeDs/PqsH
WfgmJzYRuOP3qUYuOQZVFTUVBFbQjErEVoXaAyG8C8aY1VcRE/QbTl5LnMQrfutp
B7cOq1hPEhdjiXhPspIBoIOlgQ0zZsAcOWLI0tE+NMKgiV4SvYnBDM0IVZLoHQ19
BsYXXWDOmM2a/7VvAmOryA/ft1mEwDcXPnEBiX6+FtBPKTa73nR/AqTNOgr8G5uq
PI7Aa5MzOQInRZCc+h0hdUfQ855HzrfL9ZNU2PdJzY0eJkhge6h4/WWudai7b5Ss
C8kUhqG6dwAv+6lbJZCOIcPA71VCDhu1TzkjUm2h9mPg/9aKVY0mChbh3YRkwgMq
6x66drRk8LGBKa4McxmH43gO9JbYiLc7h8mABWSiw022djPT0bxR1zrbUXcYOYDF
hJXb+MVHrhJM01yofc+jCzRgBu1Vri6F7UUW5optDH1/1WwPjn9wL6lfDHOKp9Dn
Y7zLCK/J+cmcsrKxazIW6FFjzbMFatG7Lm87MxN3TNxGUqvkekRKfHBSROGy218w
d5+uMaFWiNH3E1KJ5cxBWlQMaA0/Lsw5owGIQyqFKCvT2zAZDD1yp4Y7+KUFEn6c
7Q1949JSaCVxxjoGwiB4ey9NTyHGTTJaq0VusmOkCPqVZxC4IOWozQCaXyJUKm/y
qWMTQZXPEvGnEYtUm6TSJbZmCEFxcgDC+4hHiH2xyqDCtJY7HuERMB6i2D4AU1DU
lq1W6tJUQx85zCzBwX0DjFw7ANgZrCUzqGWa2IYw6B7z9HukOUeUiXK82/c2hTGp
yR9G9UtH7KcPbP+95B2zG910SH9xVfOfhc2v3lr4iz4wsscqZATZxVEh8R/W4+lj
/R7BJej8YMu9ZECV5Mjw922Yio3KzmZHR+v8N3L4NjyipfXywhtZoeVuZKxwv16m
R3KyDaajgFk0tGNn4aVED097W68EqWKrlAdVEL+rzmKcP1hAaPCvUdtHi5qaGHMp
s5kO72e0Xgmo7/GpAi3KoQYnc4CeF5gEpV522Akdl+gQ8FEwQbm5QNTQs5iD/GiO
OGcGk4WEPAHA9r9GzmbsePrcwGFnUCe6E4LoxshJgkNLOllhSWSPr41BWg5P5u9/
ZLmI1JBMgSXg7bSIeJvYQeqJK5V+5E0DNFQQXR5VvaN07rJf7G5yY8/8+y1qiDr3
GyIZl2ND5X5Y/nwvYl0XPSTXWk8dDPXaPX3Z+f8ejzdVLfThWcXLwl9pWxWBGB09
GDMyWss9ajaY5HyJo4RfQYgUe/FI6I4gjox4wA+v511KFDZUoUXacwUe5XBzcHnS
WcQanjz72VR09+g8DvlCZo+wnyyHQwlzMraUWzqJNzzczVSWmlZyJTevhYs7w0Gy
/+wCupQ2t/3NZEbJtE8AZUP7beGxxXldGvTnwCD5bJJMSkX1c90ar0OEi4IfjPWk
PDP6rXtiPJjV+vVISyhlWw9I+savrWdctGSGxLHJxAZjcNvxiglJyQgutP+ChMWy
qN8oJclHfnWLf+klSzXDcMuAj1MwUJyJqAq+xZy8fLglD2BFOK2xsWoKxhXYHol+
rivZ0j7vI3L5fUmgZvmmctsLMkBCA0u9GC1pjI+f65bvkC+2ox6haaldWvkV1sot
c73V+vA86FpNWlV45/Fpg5il+Q8rlEcG1w6oipsE7tfA3COMp+TuuFY3C7Kk0fjB
ucWWUMw732L5kiQ7GSjf36muZe8jFEOeYIc55vubpLipTabFbaEuibN2AB9sOwIf
JTDI5iRQUgTFBQ4RUgQ4d1pyRv/msL9p4+8FIFNHoHWx2kGEQALODezZWo7CsQo8
wiZtr27D55YuglVAukTAQCagKeS1bNYqtoyGPOYoRLU1AnGQN0HipErhugrF8p6x
c9/2iRHWhaFSNZx/fXL3aHIfPl5Z3KyhSCcv+qnJlTax8taaIa1EvlYvTBXaOnoc
At3yo0Rr1+G+9dCpv1hYiTNYMcz1CgYC+E/t67NkEBjAWfVwVTXevoiKq5TcfhZv
bjN4l+YK7btPy5dO6s8T8H/N4/LeOwNSjzZJzkm0aA4cxDYGB4hTtEyhPQvnAOA4
75zbwciMut5iRbIGtIBmS/OJn7QtKhHS6GnkDFCZV0DD4Y/frHV4nUYyRWIkLnZy
FHBdvBhiHOX4UsNxudd9ahzkCuJQqw+T7ZGIpJbSxiDit1XlEvQmML117Rhrvwol
N2tUVFUqIoyqxr8xU1VNvbUbsgE9VxRV8kVUI/6CCi83WrmNVe8DruTLtD34x70S
qVRY1rNB/Ju+BfvbuQJr+Ew2rUd/u7j0skt09ru+ly/Z8xDnTBG/Y7jci6skfDKp
L6cD1FLQYdET5yQMPYQAAqxOqd0I8R1ND4I8zXA1xWwIjNSdQCJRR/RPq6Ak13WZ
fZDXu2TsM+cGqA14QMNjzusMXbPKF9EvqK3gMYaLeWLI5NYdlalOAh0k2hzpwVDd
qRfXChqAG/QuC7ovtSgmUtjEXr1QSmTsfK4JgeSXImwM4ZdHRT0Ej/9gXD8w4E7p
45UY3+vkqGh5rLXjw4OU0FUMMP82XE0BHH+0yVfE5TJebqqo8sh3yyqojToOcGqE
HvVxuLqx0DQ1gSwAg+PZ0F1HOHNZhlETZjhJwZqejLqHtm5hdeN8OBJHZsGrC6OI
s5HwsZVDbiOuPTR1UZ0fa/4Vjd85RBFyYsaZ4J/snJTuB6mv5GySZdKe13XmRAOm
Vff+YK3UQ9xymHDdk/6tJxOhnTyHQifpdQguekTGUtyF5oVR/xV8Od8eBApxidTP
x7aJjL/wSosgfuJC5VOszUsfGrCDZ7JCHB91fb+e452jxCGXIAQE3bcjc7djPUHC
JP74R8kXCxQPRyEWc9yL/4DyTIWo6nbz6NOb1x0YDLtgCTmGEKEg4/rT9VT60IbM
ffiqwsyql9ldU7Lhjf8z7RSF6GPmUbzhih3EnAhyn3fz6LPt2obBALEYX5Yy7Nhv
fAL03MFhbOD5OQwgQxrN219JaIaedWIe0qn4BvpWEdpagAcLRJV8SxXttlqdgkAs
dHBxYTjuW3MUBNo8rAFyysWBuRkZ5Tg/2D+Uv+rcyeG55idaz6HQylF2huL/ygMf
RBxnVnTL2nTPeQZIM06XjjtrHnQUxMDYVWdDeK2LLdP/cjAXVkk7W/mO19c9fqce
COGaDFhziw8OyaMIFKfbraROED3vHyopHw/ksm1/viO4kC57TWaH/3hQpQIzKWS9
lZi9NZyvp8Zg7zxeuoox8u4caL5EgkTXgBiqj1tD3prmuErAm6xci1baiJJc7goQ
q/klSOwD1H2Klb424AbOY+/lr5Us+qQHYb1o6GcXHv3KS3QWbrmomckZQsTtyLMB
v93Jjh+VyJwOdxd2I427VNqgze9HC10WcdxUeYUwyisCYtzmcAw+QGSRsMArcE4x
Z9ykx675wLrXxFeXfGPOR5p1GGpvAc1Op3e/QxM22eD1H9ujITE7fqXp4kqIgTJ1
3zJ+0MprmruZRPQ5NCTi2dII0dbVEyB178/MR+6JhLqg7+HE3Nwm2C8AL7LeAxGV
YqRxeJmfDrL/QhnZTMoJMJU+4Y23aXOEd1gUSpQsqElq4fEyQgAU+K5GgMJVWle6
Y/fFy+qZakAh4VReT1ESmiSfbThoZoe0twsxZhhwmSkbUanCQq7xy4+N8+tjWmup
mnCnTEvMg41GF9Zr4Ur7gydRTBCgUUfOm8ujN6gZiS0EvwFMDEMifN8fLCZ94MS/
Kl3LAzGVpW/7GvukdMLXe+8jJ5Ocn85bTvv340LSKrvd3jMmVXcGNOpDT+VBI8Ia
eEn3z1Zqrzo9ad8v3ZpsJx1bHeTpQPSHMSSdGOMhZghMsmo8qA3KNaq5gLe2pw7v
OAwAAHGNtGNlJT5J/BIDOvBqqNmBep0v9aNdBUYsAMIHpSFh6BEy8uaqjxVeKyAv
GcxaO0hNnwga0jWpib0QHssb8AghGfhPD24MIB26rIY/6ZsbJoGLQXQkhB5STg27
3prhN0HP+GBut6vShXJfwiedzoUAy2OFo15yGmTXGULJd060XNIHrKg424pRhRRL
j6dw+6CJgNUm/Rk0jCeMk0Pl2rheQ8N6CH5jrkTxDlr9Bf91ePMQwa55WeyQuX1O
f5n8YhzVhf4poQJu+t18sbkZ3IXjO+XfZFaVJbOwvlhSy3cUvC5QZ3O8WQhqt9re
UqoOi2/Wsd1BU1mTGYNAPA8GFLiSlpUM77O2zlBwXuxgYSgk9lk/j/8GWSa+VeMg
lkw6WuniCkC3NBhkxqFu2rQwywsefMLj1KJQpI4J5Xcmj9PUPWCsQ9im9O9CSAfV
i19nOkMr2+OWElAUsksakcMflvdj99tTWSgcUVIjpbXfoQiy+5ZHRYazDm2ZdQ56
ABlkG5UaWJQysRAUUBBJfgV/bQ1lHKGq69g4Kpe4EKP6pXOWWw9Yx3LDnXWfK0GR
RnRT/lszMzS41FfBjbop/gwc03CczNVaTVyHY61oANC6W7ShomTkTdwzQTXm9W7U
vXRRcqSMDroXZx2IevGHfV3UP2rWOPKPu9UP77kG9CNCYMKASOzR/bT8vyGRHnwH
dr6l2GAsSspzZZTC9/Cec0bq7REZIpnMUSzTSVb3LBzFHNQj5ZkRNVVRJs5bRANR
KjD9yjCxs8cmfNfNZTBsyNxANvrIO0tPIddcXulNGxFN8RyxKbChusldfZZnOiSn
slkxOMMQyQfXLbnsVxVicDzhddKPHY/aXhx3OCf14qd76qiqZUZsvjd5CQUtmAGP
tOforX7Pjgcwzi0tlI+qX75ZG8UKo5vysy+8gx/R2uDR0XlYl+Mv/wuvMMK9KuH+
ZF/mDMYWX0L4HYGPADUec2DiEUiEpdBUk/mkVCT/mdLo4b5XEh2txFOtfVAGvCdi
QFQX4t3600klcNvOMEX/h7+y7OPmybjSSyFsqYb7Mn3F9woc4/6xvFcDzkjJeUMs
C+Izx/QyAgTgDfJrk/UvjkKjtG3vg76WC8n9wQMDiTcmwd/YjmOPiUwR7hy2JZPO
1ma8ZFHdksJ5dQ6ygJNa5bUkcZ4QnmjIUbxmlYFvTgMTJp960I2OXa+D+oeKzuLi
F/OaOLMM8Zn8tbgc3RGLl++YKhaNIIsLtIDO9vUQKlBj4WlPhtiCW5JczlEmG40u
yYdVFI4pu+c2qIl2OqUfZfZnrPoRsBFYSTj6p4F7a+eHmPVlfw/TGQLG+nZnYSHu
iiWlUhELZWZCZDV1mqzogT35ie4qrfLVI4u2uvFI6KHkreALKWcWFzpRg89KG3k1
xQ+Iq/LG/K6jMPBETTUvCBXJBe+b5tRPgEFCqvXLG5ROkfBft8iFCPb/VU8sc019
3EIC5235OsuuIt9LUusOjR6zepwqWepcyROGEOMiEX5CY+JwpueetJ9Vy23FOWYV
n+JlPegRPGiEO03ck4nYi3dWnTVsEP57vvmviCnHpZ6lYLMalBdSD6L1KjLn/852
GRuP8OCOalEXHj0jkPyZdLUt15K+Tu092DVLdYzb4JSonu7rqHsAjF1vmN014tJr
/pws0ctJtnyrtDFy1iHLgJ0ksSPTp2c9MkQNVVbUc04P3sSpdt5qIeaJkJvEsViv
fIwKF4ZeGzBtxhWkadtNZ4RYK8T62czlJq+2/30+QKtt25B6D1ZuPASokNjPHj5x
1zUH9KZPYuWZpWOrnSxi+EemHEEX/M2HTgf6ZYb9k/zq3izv1fS6X2FCSIywiYea
Qt2M2NtU2+xuO38Sqq1QzdVRL3weH0x91RjtxWDtu+R89h0a7soAaRRa+4REYiCl
U4lAJA8myHVysryCS8krnKAuZBk2/uQdrACeV3LDxhQh9JYulPgiu4zM7b/Ac7FD
nuN3EIrlbRD2VAM9WY7iQAlYBkkJ9gOi5Y8uwox9XDAgMpDh0aBYGBpetpZyf6r/
y01E1UhBDIJ3gvk6131BjIcbHuk0fOdx2k6iEW7ybTgql1l+35FKSWs9pZIDrFM3
dsxI7/jZdYYuA6TE6B7Jxws7MJI8V0GjKJy4d3cYIWxbfUtxbXOGMg6fUcaDKVjy
+D+3Rpmu04pauFDNICurT4CtBxtB8oOKZVAkpiA/xl6P+GMVcBWrb99+2x2avP+O
5CXen7VO0BAClJUNeu3Rqn6iccLrejHL/PVnkDajgbnEvU5ttNNOI5rfXtNsC/si
TjZoo6PW/6ukpNmvOq9cR7xOJSiivXFmFstrXLkesVsDGuo9xcX4MsKpSD1F8isr
5CDj24/bhG6WXZmJoIBPX7v6La3SiihiehnCG4o2Rhqtv9MPhRoH3K48EhWZ3HHP
I69k++oQ7WMHESvU4tmdt53aCO75deA0LjzgRrsU7iZ4/0AIOBXgaB4BGxxbpc0p
TzvsKZ5iYjmpOaPnl7ZMMVu8lfBVsBSSA4/XFIWOtdLQ9MWnd9RPJR7Xhqm9WC6i
O+pxaDMVB0KF0kYAVJ/xX2FwZ3ZGaxoyIIOYT1O5SHzgwpxz0YnL4/wRo4+BrUy8
ppAru86SG95pIMZn94ufiZ6ahDMXngwdpf6s90QuGDzDuLqxhInxJmZY4KA0DpAz
dXuEN66CYejJUbFl3+pPRZqJc5crwM7CxUIdngV/mAXVDExPq7nRjjZRv/o+GLZn
7p5EGUShbZ8g/af6b8xO6B3OxcZvW/2M15GK3WHbNufiRNuhayO0R7vZL2Rfz2pz
8iKkTwtQMhzyrp2P/t19rJWCBe1Rbb2QNP2l/OD3vZ9jP0E/H9ayrBLw4rK68cvp
fOC6l6KbfbPSpSL1Ck+c3mydXFEFZTEvHrY937FSs/hopdtWpByoQpDig+HV0Wn3
XpMj25W/itXC8MUEXBE0rPBiHoRll2nuNsFvZ3nbTLHel2vXrNnJExQd6C81vtOO
1uhYhRnMFLu3TFATXCnENBred9QL69YwybYdbR0AZhKGb9npPXQqLXRvvy4/3KuU
8uImCE8i8OLhRWCTWQgeo9AyvV99ZNv4SUZngO0pGqbn5m+oQUHeSRxzUAC9DNp8
2LEEKLrJ3Dxu36wvMPZlmk5h7qq4iMbmMUu1exT3whXwAyUb9X5JM9C72qQ9Ha11
7OvjLNUVNKu57UBaMVuXwUmUH2z495FQfa0qm1s4ToZr438ckTmequC5Vf76bdw2
+/oLrRKE3RpQtfjmM9ZItnYWfCGCNvbDzn24Mi1J8UyMOlk7OQkwzf+a9qmk9hr7
uIzXg494p+p1eek+qPbmTJHgIgNvlZu5q1SbICjY8LXBaWhNLWBkvIjNTR0wQajF
Ea6X4NfRHY9/k5tp2f7c6bptKz4rPl38lYoez8MOHXQIDzl20m9wg8QDLYiBzgMe
gZ/g+A/dNQSYW7sF2ohtoXectX27y+950HCNimteHYRFBnPG7Wt/OzZb1B7oJ9F9
8dMoQEKsjIAUIAs0UsTM1MSR0D4kETcgGsZl98oxdplrbTeUqX7hWCqDNAaMpTjq
oZN+BWo/9bqaSPcwshO4turOCxuRzaCJRQu/huT8JfC8rxSpADNZ4pOfpCmTnMRu
taLJaogfX0ESmrgmG67KTHKZsa/h0fIzKafdJPECcCNq+tM3c8IYsd7skdLP51TZ
ahhlSkEwcGEPvJjmgNYOtM8fOLbyIwYG3+L1NLfBkp5d5BNVBO+MaX3+LsNzPWOK
aG+Y+gCBZVsxnHDnEKs8ajzTn81FI9yQF7VmOdxSqnANZzV15duzyZ40kcmn5D10
WJMK/TrIzYy6pyRB1ctDJtzH3R8QclO1zcEQezlbHG9stiaOM0iyqsN/tbQMPHts
UaWPOz0bprwTmafUX5jFynXK6WWgjK8aFszLyb4KHBaI6x81Ee+dOt1aUFVIskW3
k+sBXmj//ocxW0bjCM7qF/vLyBJMGAb2GtuQdZeqStzxYKJtOASzj1Y9heFK+Pj6
heLF4tw4ADtwpCqdsveIvpkk/BHukGzSz6de8+Yq7/XSgLXeYPBkWt46jbTlzhlL
RKQkZRu4lrR5IUdlfntyE2e6/rCt1tZOhQD8HU/PY7O9irqQBByu0ik/XZiVJQYE
8Zmm4pO33VHzkmuOp91G32oZrbPpKUVX5kfte7Nu4sv9O26XOXC3eZxEJOifN30P
RqM92flRNhCuB84tT0mMogbsrhNDK5cUEdB88XkwIn9Qe+//yAohjo/eUdf+4/7g
MpzqkZecnL91iayxmo361Gkd3wOCeHymrMJ0hyl14y2tkS5lpX7jRPCqPRGG+esT
6WCNk2VzU7hQ8Pb/0R+egGGH6Y5+83XWmCpaYAFCDtL/mV9EB0OmTJNU8jj8Ss+x
6AnYrq11nxZe8o7GtWfjjd67LTi0yjUIHlSoeIigPX+vNjhH7avTnIqEVpZz0mQF
0GEJexHj8YmYyAvgptoqfVc7Wm4zdOJ7GmDZUhppRbV9OyqsoXOnJVl/OgNwK8OM
eGA6le2moo1woNDJJXCYzQzy0FoY0y2K/3bQ4+HoLIHTSycuhxySfxoi2OHXZHAn
LC40mBIlkdZFRlQYjXhWQwGgOFBHrqzpi327jLzBQgVyLj6cUCsGL0T0mmBokvOJ
SLqsTEYDZ9tjTGiU3Dt8fHk3/rb2Uw01pPMS4b/4s1ejIkSly7D5x5s28gjd2W9f
E2YDEfc80ZyKJe9QKTdb1lH5ga8r7hdUul03cO0brWuEzT7mhDj23But3q5oJwre
lMQQxGBM6o7XONRyf5LYkJ9epNbGLZ413aYT6pzpo29+j4C0C3QFENJ2JaqO6JI1
nwb+cntjhI9m/ny213RsklxPdk2FiLpysIIWNhP0HWEjRZE9f/E4r4VPVdmwUWMi
fZoOJ49+jELBsIpFD6M/ZH0HUf9uG74dPaytru1w356hRT5Dg+bCuZFD9LeeMMZS
pg3U+z/a1QEPRTDzjn75gqW3QZSmoana0XNlU3QAyH0V4H9oT2ghnkoo3/ApiujJ
4ShkDwdqsc2qSShR7PvjewN0eIHfnUuDcpwYMKkw0GcoTlDGktpridNDyt5N6rN4
yVyNnjOXpra+uewTmBvN3U4aFuVUS78F4R9paGONDEx20bBbya+vsobNSK0WIgeg
G2TwAFVWKYsO3tObKG0oLJ2w/jKM8RmxNrj0QgjbQkeJ7MZW8OFwX7MHs6H/x9DM
qeRY1fa+dFjTDFPhdJJERfdJTB5UUCaPywzE88UmeZWLBMb/bfU8Lcpaj0k0KKGo
/oO6t8d/F5bo162DQRa2qhcVfYsADia7dfSGS9sFgbX+Abn5b+IGZfhJjt4Pl8YY
F1kZt/c7KzaEnitJWT5i+9ykhWPN9yP05MkMTaMVmfTE3YVWWk/HnyGFyKgaBOIY
WUn1wx4RSpQ/FWaJuMjPC2meMBzdaDW5zlQjsWwkcXVmmOR37lNK+bzuaXoO7ggO
rNFOsAz07oX7GdjIAZ51ndSBHFQiBCjDLwWw5KZV45uSdmczQhGhUCYP9VqZHToh
hmWBwFCHJDoIlTa/tV4FDzdHhuxG9OMtsq4CeWPQa7mPMq6Uk0Bo0T9EiuXROtiv
QhB8UcgGLd/OE0HiIUzIHL5guTnEKJkX236vdkDEG1ZewphSHq2xJ695Bkero/0F
boF3FPZk0UJ/bKGZZqU/y7HuWCQ3RXZs0MCyhGlHyR4LPT08WdYbboaAW1cNEw/j
C/jpOB1yhumpsWtbBm9Wff+78gNTk2Fvv+qSlX4d+xHTe8DBQCtAPqLU6xsQf0s1
LMJ24SzpaosaH2RpmT49s/LBBkR6WoicZHfgYbikk0CxU/QilSbbpfDF1sEYfSrY
a3jYgPCUvby97FrWhim5Cmp08W6zzr2ydfcQ1hH6x9oiO6E8huAVARFJPTSLBcg5
zZGgAD3Ygxn7Vh+2wUGH2DsBmyHawaCEZN3xn5FQs5j+1f3u2wNta1JISXpgEI13
UJDlnqkzYY6fr0wirs0ljw3gznr8DnaPaPpjtqvWqe4UarOzDfHQamimJRkuDsDv
GGWn3P4gNsrexYaYCaZNjsVg+Sm2HuCNr6NI10MjGDAbwMkFr7XZRr9cT6K4ek8Y
ix4Q7PP20sq9ar3+SJmo2wT8kQGo5n5U+juaqJFggV/XGo/EQgnR98xtcKmWO6j4
kL/YlVg+P0rSe01+cnYC2uWHZYuEVoQwDDv89a1mDvEry+JFnPaA/il4va7BuSWm
Wc4T8bIgS5QvpdA3QZaZhdRwn2BL5OaNyNIuDoqHbDWqaAQ0uF1YUl7b/fBWX2/U
okcxy/3tWjsedw8O2JvsWit4Zme/Hh5WaBdhNz9qdo//cNvWxFcuIxnDZPmY9oqc
wk4W30eaVTPxtRwDwwEVb6o4VKKL7kcmIhijdzkRArwAodl8n+wjyDByFYPCp8Z4
TRYYc1mGuqh4e/kVJ55fXSm5oUNAwzbeKAhOUldIHw1GlOrw/c4/YJamADQm/yhq
/l3szO5UjKq0L5SoIbN6SeHzdUNJUNBfNkyYkeiDTzZAvV6XD12RDv/WX6kTeXeU
xu6Cw4f/w2ybfC9b/S/D87jbgqqYQUy9BDsAyfBIejr6Mn1fSAE3yZyHBwLlB5FI
DbazsdbRE7xs19LvcLJywyP5ZHm/pYkgDpR1720JWCHLRtjbg1TobOKjWhLoNW8p
8C54fZCVOff1lPcDxeJYii5A6x6O9V+2wZK+nCpsxcwapsmSXaybbtmMzM/MgrcA
+D736qVirm/B2rF14OfMU2NS6hXn/IuD13gPrpgYM8BeFBYxpZYoO8sBmmHJg70p
xE4zs5tVPV/VNai7ZILymKBMHjqXNHX6XUhwgFlKNLAm+vWioe23SMLarrTrvy5F
hImtEdmXcpC/lDSW+FdYOmyY2KcD7Nc3PfSfAMhyN8kMSqIf5ra8Xx4JPRIwnHgC
JBE9KFXstZVqUQFjHIluEwfX6zZyZ1yEzeqWU1LNr7VhONYUbRwQtmmtoQNysipc
T0AOyewdiJNLqHjx3EdaoXQiWfdkdugT4wQqXQwxCJHxPDACfbkPVuf9sVsqBOrU
Fg5yYybrY/DgoaLjRo2GsA==
`pragma protect end_protected
	pa_bus_tracer  #(
        .DATA_WIDTH     (256),
        .MAX_PKT_SIZE   (32),
        .PROTOCOL_ID (PROT_ID_CAN2)
    ) pa_pkt_tracer (
        .i_clk              (ref_clk),
        .i_rstn             (ref_rstn),
        .i_header           (frame_type),
        .i_start            (r_frame_rdy),
        .i_end              (r_frame_rdy),
        .i_valid            (r_frame_rdy),
        .i_be               ('hffffffff),
        .i_data             ({pa_pkt}),      
        .io_connect         (pa_c_handler),
        
        .o_frame            (),
        .o_fifo_full        (),
        .o_fifo_xfer        (),
        .o_fifo_ptr         ()
    ); 
	
 endmodule
 
 
`pragma protect begin_protected
`pragma protect author = "MED"
`pragma protect author_info = "VirtuaLAB"
`pragma protect encrypt_agent = "RTLC VELOCE", encrypt_agent_info = "1.5"
`pragma protect key_keyowner = "Mentor Graphics Corporation"
`pragma protect key_keyname =  "MGC-VERIF-SIM-RSA-1"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype =  "base64")
`pragma protect key_block
hzxUyK00R7rDJ2kWSJjSmMVTNd+kQAI2H7i/pIufEaW8Ah9RfJQoYEBSqf/Mr9Zy
s3eYTniUkNUpHGzxqAUzWUpQ7BrmLXI8DzT+NjAP2fjAvP4+UdZV/flgxGnmYd2I
OfCdrk/4V6HaItq8G/KYbFkTtIC7QudSENPdmN7Ze28=
`pragma protect key_keyowner = "Mentor Graphics Corporation"
`pragma protect key_keyname =  "MGC-VELOCE-RSA"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype =  "base64")
`pragma protect key_block
RLcX8g5CqLT17VwLeV1Y9SIgsy1Rq9DZ6GhX8FA9olBqOgDJWRA7AMzgBL/ABy2x
4iUDMY9GCoQ2otjV8G6DYpdTHePt786m6FKkvlXV8hZOtYfI7bSQ5QAk7WtpUDNE
Gme01cEiO6n1JORThKtRIn5kFt1ass1ZMhyijcvZqWo=
`pragma protect data_method =  "aes128-cbc"
`pragma protect encoding = ( enctype =  "base64" )
`pragma protect data_block
woYd1v7s95eQN1erCNe6Pr2fGIvJwA4a5gaaCTHd8IqA29m40fXXGXtfOeWowTCS
tNhN4i3iuaa7kUOcFE87yVYdmtzK7a8qAYDFQPCag+3uM9g1Ac/jLPgi+cWyLGw9
fMyzsDgVblh51JGQmTt1roEpFZKTyCml/N2g+ipGoKcccvrfX5HlEZYw/SRLq5B3
mZLM0teuvoYTJN1CLGoSt60BSmvXlA8UppJ1C1fQBaM9gHGr/sYz19Z/qNZrqjlp
Kj0bYYvgvhLto7njiH6/7sVOqVfvHaXr3BxJQAUhW+sf0ROQUeC4EXn7HDJoc6ci
znzIdcrI2p+/JScVKcr7658pNFtgSgVbBPn8+jTNhmhW/7isDTbbqB+6xHh1Zkym
mkukCoqTOjLtuO93FYljJ5mBWg2MisJ4c0zJ0EByOBP+WQyo4YBusF6NMJ8c343G
TUe/2rBf0CwmTRVYRYLM2F+sySx5FfVDeJ5eWNN/6g+C2EIQiHk1pTuUQ7SjmNSZ
KmLmcWMP2lSk7ss/I7wqMMuwICANiNzF2pDWzb97RLxbOS7Za8ujfyXsX0EdaH5s
/T22RuAVounJXfGEvlqrtEiZKKipfTDCOubZmbq4FlKHEqC+8nJAXFFzfa7rX+HP
o6Zaz5RUzdOtWOplC15OmeJ/iYK8tUEs4ztXMddXo+L3nNseUu+2nqAS278qMPQg
soHuVurzGRNlw8PXm6DuKXIjiiM9V9SodWUbkZsAKUQll1ObXBzy5LpdcvW8vurq
kBsLluFT2wWUPNa8ngCw6zcOPBML9ymRqZom5rgRVsePaLvxCB3wrsgnnRFKrnpi
WseD/zcQVG95BcQqBopwQ0iYQD0jokOA2nM/wuT9LXyQTwSlbylP/TmLUMkX1nNK
8tRugae31nL1pmCe1Poc0E/GjItwFt1+81qsmUsHVG0rzkfYmv9G1LjqSqbTuT5W
eQUoWv/bwiCQINyMq+W72qhz2i4GlWZPA+3famjJqdu8/jI5/LFstCDN+1t3VliE
Nb+ulpfDxI2hzQJSjwrf0Y000P5BOOe571xzMCoC3QcdHBjfu3QbY/enJIRiDTD9
GqH6NL3JQG4fz1EXOm6+VR+V0j+Fd1iRLSJgPUXdkvK3T84J1MWOaYiXu/aqvhLM
7viYpayPi5G10BaftiOq5AhmI7P5sBs5yhAThOW3nnnRQK3d2FUVvUm/Lu688LyX
hPL8Aiwo5U3xRI3GlVtrWHQ7OiVKm7l48xh9UCm1Jq3a+yEmL5r6UD3zqhRVw+y0
cN12+ORbjfIftdba40Cu5nEHUfZcpXdpreUWeUr3ysmyDqZyetmavlze7FIHaeU8
tysOGhALkdQvFIhrFLAzkaJbELqkwIjjiH4mcZMhfQbM+QyQYzANgsr6mRj47EBu
lrF54/YF2yLoapJPIePvebdCnivqhziiTpoFIKdz9vDY6fFAjTWFFuXcIR/6fT3m
1gtpcAm1jhCVs4Q7B46a0QWJYy3mMVrk+j/q2gj9kaR2gusiVtqq7aAcDSbXJPSJ
7DjSFob+7urX9sEYaLq53w8vCKxighmk8bJUjHCyc087dwwFpKfZVVU6yjKITatx
9LplTw29TT4RSEx0lE/aTymFkWpRUliPwxfXQdlmRaqZV8KcIu3dg4bWOexKq89l
OLVwfOIKRX9W3ESHEqtFh2vReGD9UyIrsrcYa1UXtTNnQnIBtR8uJHa1L9VcCvv3
dv2T+cqE1sE+Wo3mEXdTgLzY2R8yhRxxdpJIN8DqA1eLHauXuxOe4hlWnFrtv6lR
+cJpAFeGn8WIZ/+eV8vC25YxdyN9/zrOsB9yv8QkEn/UJpATY7JpqzPlxZAmmBR5
97WKNpCbOacHtK2jg5oUXbT62O5H3W8X3KGC0W1NKdmdufEPAAHzfqTQe3lqa3xn
gSZw9Q5mQAJ9oZP3mwDQz4/mCrDquWkVwTCO2xlSufShifHyjzAZyUyDeKNn7w9P
L1VS87Il9Pa3mdtIPOAX+JkjGMLbVRzLj15olwCriXsG3SK5PZdPG2KL0bgd372J
Zl8IC1onI3EnMNUg6cPKR0idToOTCGK4hnrs8SA8cDNe49xPC6mJiXFtyG+iz66L
PoWmSKNrzeOyyw4QGblu9UXnvrD0wc6J285IgZBrPC3OE2m4EsUP3SCVzqrfYCpi
6hAiFJIfoxCITz7u1Q5nXD2YlgjRR9rnuPJjTUjDJ+SMHh/m08MqEQrXVSAlMgJY
i9hk6ryVRo8DOmoRUt7Smt8YOkVHyj3gq3a42fT1REK3oYr9c6FMRwv4raLGLyxv
uU36XZ4vsgWOZbEf12/MNE+Ax+npI6uZI0mWr5LUWYNJJP0EraevKEEE/53zeEBR
VmY8OC0ZvUkR/FqEQaIxOx7jcoi/aIhmGkSUPzKA9YZXGh3nM37moCU4SJeWRy+t
BYVm6BjTykdK7rPyXvWHZrOfkfwvDA8xhScRXuFuvFegIlHTnfR6FPNbgqmbH258
cCmNStED5cUWZ5EOgGEIVWtgDi/+oWMRK02Qswy6IRWPtluo8JRm+PDrH48V+NJm
w6yr8NYEbdGC95UGFJJixo7VdJLRjr9EuGt+AAy5x7CDvuofOGIs5M1kZ/hSm+IM
8eSsGqssrd23vcg4c0JId4mTItsAk3kbExpJ4cz2C+MfNIVCdLojNqecUNdEBJ7n
UjFOyQI8cw7c6ylnXhys2qoimfvonpXuHmbQugWushGPdkkNHoiKVm0pHrzHxsSb
SloAgSAWmax12llJNSZDyZldd3qD9eaPGUvJR+UPteZOr0p5F+bcwUnd1WJ4jL82
BaHMmdkbP2cH+rT/0jpg6qTu3n5wop2swyQj+3cGqNRpAOONgP5gl//SsrcvJa6E
nQyBiqgoHNcFkjYb7h8JUClHGLoW0L8RZ2CnpvaIWTH6vdWDz8QmfnK/GnouNyFQ
rnkh+fTEs1n4lmFIPxAauWrZEeLxzq/caOImIdkxrBPvwvMwoHmVyjIYO/lcMtW8
vN2ZHLrWa7J3olegPYYSOALHnTGD2yOe7tzF9sSgCWkwFy5ybnjtOgpmB/SyID17
Oskx/zLVW09z8A2RfvsKmUSuJTs0vUtk30Sw6iuT5H8OEUpN7B/tWZQdQXcZD7Kx
l9vVHes3KGgT/QWQACzB4f4NPWuk6xvZMQPSVWFNeRb/hJS/z7MWXFqrNdZxwGoq
gIETxmQTima93vnynVBzt+RBqR3b3OLdb+pXgSfajmXa8Z8XXaXU36J4PPMr2mYv
/4mzgDRRZxp+p4x8BG1rZiHhmLt3kDkoVyd9YU19YqwHyG88zs/aBnHm3Bx8Jz5Q
f0ZwZjcZPa60y1lALG9y8UZfTlmJMVMnNlOVwdxNOvitA9aDObr6ysUYARMRs7X+
t6C3ALbknRE0OSq8CLhY0cAzvizVK/WjQUKGY4usDlHI1yYduWlmWwuQwTqNP8CM
RSba5zMqIixtUU860+iAc5QUZYQ7m8rX6S7Q8Z45Vcftd3WpHI6Ak3I70sMc01zZ
qwjhGjErYBs2zRuedAnLC5prtINXbid/ELSJM2eT+EKghPFTNvtBo1z/W0HS38Ss
Nc5qOYrKNGvdOPhBsNv2u4ff9pQyJi0GoZ34OE9ZfAKeg77nD+ujkdhmfq5eolkq
mNHouhwFaRKdyZ4ujvRFXyOs36nRDlErh6CvZO9QDqeY04yW8EJnrgE5gBBhIWsK
VsjK0UptbTteBRdtprV4T+bbwBmUKVUlWEf8JH/yNGlVYwt9MfmlULhzC+65JIBc
Pgn7Pw2asMbXYjhXRU8RL52ywsM7lv3oG+AaawIQedp543uTgkDOZ5c6GH47/xXW
J38QR4+8r8hpPrxY65v0MGe0DEmdhXNxAPXJM8jU9XDmHS737rOG9Gq6WXVY6eY2
Bna+vAtES2o/ySoH6Z0/g2G+fXfvt1BvltVGK9f6XxdtdZxHEhF9HlGxtzQjdIuT
SwRmOvuf0taSlhKIQgcEioWA3aj1CHUgJqMqXzRBP2Qxs61yKAB7+1H9Zjz+v7o7
JLiXCA53avaEI28+DA+RfJzV6p1Ld2SYEPX//xwxSfv46Wfk4V+jrwMuQ1f4VUzW
15XzzqctF+cXbqo04Zz2Yi1KCGNwWMcO2mHpN/fERejWKC47aEc37UnX1ww80K43
swk7c0xujEaLCfV58zYLuux7JXpirX0qfKSKqKeLDZNSPmx046YuHHoj4FHTKYsH
LeiTv1oGeRzcl1u/rbl89nFEMT8O5RMNwJ0XCn8edAi5AoEVs4yBYqkm926iGioD
WyuDmXPCIFEI+kewFPuLzg9jkaDVEBUjLDKtYt9lPAktsC8HZcvjVukyH/z8qm0H
`pragma protect end_protected
    /******************************************************************************
    * DPI Import/Export
    ******************************************************************************/
    import "DPI-C" pure function void on_pa_ref();
    import "DPI-C" pure function void on_pa_rst(input bit [255:0] param);
    import "DPI-C" context function void on_pa_session_info(input bit [511:0] info,output bit [63:0] dummy);
    import "DPI-C" context function void on_pa_get_chandle(output bit [63:0] connect);
    import "DPI-C" pure function void on_pa_set_chandle(input bit [63:0] connect);
    import "DPI-C" pure function void on_pa_fifo_flush(input bit [7:0] data [0:BYTES_COUNT-1],
                                                       input bit [31:0] bytes,
                                                       input bit [31:0] pkt_header);
`pragma protect begin_protected
`pragma protect author = "MED"
`pragma protect author_info = "VirtuaLAB"
`pragma protect encrypt_agent = "RTLC VELOCE", encrypt_agent_info = "1.5"
`pragma protect key_keyowner = "Mentor Graphics Corporation"
`pragma protect key_keyname =  "MGC-VERIF-SIM-RSA-1"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype =  "base64")
`pragma protect key_block
j+L/WpLxyl9wl5h4ErMsUgGksDgBEngQijXBqc6ooZfejDfsCaIZRCHv9JEyG8Wd
8aU1AA70szirAS6IimxFAv4gDdCJdQKt9Z1GKKRY8QKQIb9LKFdEA0Og8YYIXIZ1
PKYpFQ9q/XXyI9Wnp+8isYQEHRy3FJsnBttwC68oKFs=
`pragma protect key_keyowner = "Mentor Graphics Corporation"
`pragma protect key_keyname =  "MGC-VELOCE-RSA"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype =  "base64")
`pragma protect key_block
WjegJ4Ewza9XPPyxqCjgWxQFcvg6zq1Plp23ISh9W61GK1T90+daY66KPecOGij1
Pv/DR0awHFfveyWWZ+L5MHnvu3TpAAJmhqovyvMhDeUqCtuKIbmQ4Em0dChYRfIl
8GdiiL3b887v6TTWhKNU0zjSHDXNdVNSyvnbx5uWQXo=
`pragma protect data_method =  "aes128-cbc"
`pragma protect encoding = ( enctype =  "base64" )
`pragma protect data_block
zuA5QKbez38ATIUJr3Tpe8hhW1CA22U7eBSa0f7IQ6gOIBcGjpMGBnP/I6qNGWmG
T1vjFNoGYvNsE7nd1HDABiaO5Ju9nUVKuYdZfHs38J4YTvMBFxB5nR3tfFpAabN3
+h04J5IEeg0pNkrJz7qfAULLAjE+Aecgv6rxIKH+su2F43lh/z/sUHGHUp3C9Exz
uOPoxhrbv6V176oHkagjDktc/7UMCLco25v+XeHrW++LW5VvegctyhJ2tzSYyj7n
J7c1g0+vOAPjc2vdkDv6Ees89VFU1FJpBWlPBykH26LOaiu9/VDjalTfibTlOh5l
umUvSWwHHNAFxpcEDq/T8aRXq+TqmiR84A3egGkMJeOBod1fHwT6F+FZvNA47dGm
LDbTpPxYKxLsTpIaILliCRw8powuhqMPyJEXhVfl6KAwUpKEWkMvB7ghEnlFZGmD
cOWm0zEQ/xi98TUnkY7/bDUzuvAVz2DwrKCYyUyDo0j55gqZnrguQoCV8Ju+2qB+
MSAFkuLsu+idSk3LlTkBLoPrL4V9bNg+1nd9B/PQwSJNocMoyhGW0sR5lwbGsavl
1zqkyUxHmpeuSazy+usfiH9HnQIEXYlvOmJqpMmmTxZWmWtHjuTOUAk3p1ydUHjl
AoTDwXirBHl16Z8SfdGAdhFSssXoGehfHQaSjKsmPgB2PnJdaF6m5568VQVMtox4
jhoDd8p0YoAEg/EpkVnhSpLrv28sZhQhzDIuL0gW5VYDHRfF2GP73cRAXF+qJxNX
PxfTTIzORBPBNPaxMCG9y8YLPrJO6MIg/R7yqLsten2iGpgVZy5lKLl04CX1FYrt
zXBtMUQ35lgoyde9pBwEJ2UEhth2TUFgqYRDolsavTFxgFtMaXs/ArkUWoVJasR/
y4ITr9Bb1LlQTLTRu5fB8s/KChJWtK424nElprKpSjUR/wSlGQGICx8R+AjjSgcv
fTs37KzlxX+WzKxHmfFKQ2J1MnT6Y3uRv13zDZXSqztngPYN8nZPoYQDbbc90tO0
CXU17s0BGIJFyuDhYt2Gyj9sS1G+71w18QtuhcGWVjW+4ACtNRpfnN7HPjB+BzXN
lueizhBn73sRDoo1irOV7aRONqMfxHMsym3XERY1AwgJUlqJSX15e7Z3GdxUJN8Z
A922JvKybxJOsD5pQB/JdOBP1WLJMqMkaJV7sywJ9R2dMUsIvLnExlLIqca7gfRH
DVlm/4VW3u6yLNTUyWg1sJO2B5PE4OQQYGmDOoIv0ywS4leYNSC6Z6EuUoWEoCHs
sgeBo9Yu4rQ1hXSKhj8aH80i6/yggObjOznHxVDAn5VtJJmVdV3r0PWY2d9J8p5E
yM5r9zSnG9H07WLYbGjeDbI0ZNnH+70ibQAfn3816amBjdB7eWlC2kHqlxXPA9eB
Vx/wn3fF17dGoNJvsKdoDyy/+C6LuxaTZOgDXsG9mmUzBhLHT8HMlsVzy8Q1N/6r
YSzCCk6uNq1CoeytFHWo6bXOFdCfOEujICQbOsXAouPzxCL1cVcictlsVNvM/arJ
KDz/LhGOjLGe7wu94AWDUyf3INACNDyZRgq0gyCarJEZ3WOUdb+mxxP4r5XFQEz4
vrPGfSCm+VRSGGhFI4eRWOEbcVYpYAM6lPrGkIAtoJGdI0Y3fYeCIz5d7oOdq5xj
dSfkTrSreQPGbL8abscfxOpCUScFMnbBkfaTv2LH0EDjYbAV99ZD/VtaJePtc8a0
S6A5QtyaM9if2L2VMNttk1k6hq28w00hpGVAR5gfF5oKZ71gK4I33CpCeC0h2jtn
JdIez20QrawqGbjkYSEc0RafWBn656rM6Vk2Jf2IKguMWJh0zevBBOiNMz6t00Nx
ffUscZMcYs7FJsOIOoQwTRzaL0YmhVp0H/cX/f0lES24HyB/8cgYlr2mTkSTzXoG
Rf3IKqrwCXgLCZEAMlLCNd7hS5WZnBxYiH9az6OdyieYA5RDFruyr8PnnC7ZM2qf
aZNKDHIeuZaknIt40IeSon4KzUDDL+vEAUJLurUvz5de6k5FmjdQOHu0v17CXKZE
lXo3KUttZuDEi5AD/i4Lm94s1+SHM+HZvidpebWurRljMN4kpp+gRqroVmvLxAQH
mhMmitxU1Vzl9+IGABYDPjEODaJo+Wiwxs5l0TnhzaYNDvf60/2JgFsJ9CVNwgpA
Umhpo1xdXrLNF3LmMuZMzSIiA6cOo8zAAuyxnv6We48jMX3f7op4LdUdemcaAKNF
feT92bRD2cJwCuu+gk2XeSbEo4pEkuvRlzZcEO/8a/kQhDe0Vhr/av4UCTye5zaM
Ma6QHQqOoZlvMCX4z7jvH2fonKf5rYZAXt/DgQ/azEhuD2fhDa+dahrVo1ek4RVh
S6edgKQeH/wOhRRBpHwRZCkhHYFq6CvUQMfU1Zfyhy/HaDA23/3Eu4UivyyXwXws
Lo1nhh3y9cqlVUsnesRGwmIAVfCNv31e8uUUhH5lLfPZFE99RYvwGcvRBL0lz4lB
2/weWYC8Z3TiBCABl1wADDlmparbOw+rd7dP7YhPvNHZ6p2bspn5uWIpFGl33g7I
my056ntJHwb/8dwTY6XyOcytZ+nZ0+hVTTQzHCTAvrhp8uBr94Brfh2gTqgsVb5H
NtHfp6CSIGy991zLYGs1OuGQi2wdkprFABW2kTHtFQk1YvImlGU3Ihn39w3sqHqL
DjlpkpXi/wKurgsBMZiad8W5ZUOGVI77lx1GK+exihqjkotGzHLAw4REeuDO4ydY
KYa9WLB3o3gjq/pd4HMWa4jp/rAJbg1hwdBWaK10STJOKnvc7r0zNoRC/3NlFqiO
xiPOgDBPbXIdv7Oa86rEdScb6gSOYtuFwGspPz+WPRfApOCm0mWLTm85HEOIeonv
sSyZRNeRqCHMmNE8gpXcYpTKDRHWvBP2blKGCganIUU105iRs3hNb+HH/m/DTBMJ
h9mDL3TxTFA8ogzeMFx8dbOQkmvpj5lPOFGDsMQsaKRvNGqREG6hAEq/3vVuw8Ei
YsyiV2axA16rhchy5aZoi5NPlqn6zShiYFQDT2teafnoYA58QEIstadMVwO6nji9
QUpz3N2HHmIn6S2hPDlB8QYDDqSlvVF5vS5n87aSlSNrz9KK2XES668RrPGrFNrM
qiBsDTrpCADE2j0qctA/8P3uuAGwXmXQniyHB1P901a7edbZ+JcxcAsmi8RsKQ/E
pPpBfmRvXnyFXK0Tv7+R9aT/NmW8LNh7EYeaLSJpLbtlM3n+rpWRr0RVSijyiLnO
elM08L3Osg800LboD8QGn7zslkWDB60I7NrXVtNzGSUPpby3cBZ0crj80CO0fxwJ
AbT+jymkFLv7wE3HAoYeof0YE7qhA927vbc8cB8FmM44KBtFOEFixcDhyHjYEgQv
URZpjJzI5We0sLyKDveo1PHj2H+UPfJq0vo3mK3R7G6i6QzoV2YDuJo+wdp+WWeP
wnyaVkUhdzFq5vITqCuRFq3MWbEnVIV3Dm5mWTr+eYND5lwL6e8u/WSShCkjd4eE
/HAkuy5urJk5dlFB9lac8UcVcom40pDI+BeF37e6Hicl3Oemx6Ookex0buR4h1Dp
c+WowzHxq4NYsi+Z0+K+RWVm6cPe1BpOjTouj4gZ9ZfBaWq9VT8ZyN1dKC7uWGTL
8Q0i5ygoYiQq32lZW3hEtV7NWoO01222Oa9Ft3fV2A4+xsZ6kbn8yjz69fsHl6r0
v86iL1BjRLTVoGI00E0AKzfx4JTqhSYgeyDBTJirKQYioQqIsozctukl9Y4XEs/u
KwnWiR7KTqlDRk7zZwMmmK7/iDnat1VE3Ttm1DP9+h/NVbl7suf10EsAz8luHxXa
1vv4BWab8Mgt4SNcQPRrTsf7UA2IOa2pf/46pgUSjpNiC3q6XrhchLIszpuS2HYW
3rftLMuwcxDRpVyZICRWEbHXYvGO3AlIlfTdMH/YtmCvH79sRd2UTepskbOzi+aU
YRMSghDm9WmHyssbkc9FWdXae3PP3jrXT/0e4gKKav/A6EyzVWSw21cUdzJkRJ3u
i/CfJrjy2SrEttsNb7IG4pObSbV4uTIPy7P/XehCmXzg4uULnw7qikkE6NkVg7up
dhSH9O1lapvZIiMPNSS0+a0OE4TYsL/WJGzJKsw4t53oSusQF2LEYxbuzTwms2oj
CvFoX+7zAXJ4eW9YxDvXz2hL/dCGKk9lDd0W1vAm2op8q0MVnJ1FgdRgTSMhZnis
qpTni5mhbbwP6P3vGKHGTQ22rk8ciN2Up2swxE8JniBWk/iGOZXjba8JkHrIdRka
kUkZjBvKu41nBG0CzPAFZD6eONzRFFWVui1PEfTVaAWMAF4Ev4LoeLRIVte7X1+Z
ZSpprD4o+fymZ7gB50M3WFgA5ieKoozPE0bc0dJlZREfiUPtr0vzqgDFkO+tl7fp
ug6uIcoEQZpSXkwIYYP2ugzysKQzF9SiUse1C9+fy5lJPm3oP5I2CHedwZZ6F+qU
R0mhpp3RgkNxTowYz4Xsu3wYv4lAJ2K7O+Bhc/R1TkWQE0nH/OMEeA0Ll9/njOxr
BfWvagtYexYbkFIS+Qt6uwfK1Q/R592mYZiCDfZgMHK2iXCTVpttpgyOVko3T/o9
Fzi3kssLwPRWs1jBZ24gBEvTyQArDsQv5F2NiberDLb9+fbR/OZYtSsKG6KpNsuU
ENr4tz6aTCTzJxA8tVsDQehZ/amNpaQz1uHFHiu52kfTLNj9h92m7xu8kb4cUluj
OJ0iWy00VzAtfnRD+XA6qD0HJUK6MmDtddG3MeVTI/l7oX07B3TLLIsPm6IrqxVj
qgTP9+b/SYE3kY6Ke4zvsuBnpKE1eG4VL3iIgLeDyoviGNlFvgvprdVs1U6yhXZw
jGc2+0i9H+GhCWKz6ejAg43h11OLw3/gWvxDEfYNux+sMB0zuWQhdHzQeyWnmkKa
HigEaCH8tF0FdPGF0lVcrKs0R5pk38xSAkpwtH4k1tS0tJWYw3/fMQdNfCaPed92
DdmZ/lDNewqmeCT9Nxat7lgXwbyPh8Mk3rhwD716s6oEE1kYnt3hXHA7DRuANSYd
wKTRx/omu4EzTsfQ8PIhc+xD38Y+JkQP434TkshF8uzXlX4FtDRrejRgdKnyQYLs
HSuHTY0NqCiFnMiJfTGcHILJ+rlBoqsMG/4awBI53dhYLVS13UUFOQFCMEyZJTio
4m6GxVxz7j/0nXvQanUTlo4Jfi38t7C1Hnc/t0u3q6nAAZ7F5XDvtcW4wCQs3HI0
FlPAuJcN/0bN005Xh4fKUbVI3BE5kezPW619rHN883bXkBYB6ierTGGNDeZ2sEb/
vHEIrJp7BzQlUtt9uFfBxSxwLG7Z8RqPxN69Txw0LW7rotnU80iy+Dt7k6JMKl2J
SrImjxmVBVTadGtpZRDnCncFDOCNEYvah+5TSF7Vc6bZGn/trBnxhQfBbH0QdOVm
4VEVuVTpMZtU/MdKHTLoxmWWwAgmcPe++aTxODAS0Ds5CmoJZ5WhQhoZsyfCueis
jVGinZOBUjdTRdqiBJBkr825xENTFyYG/dsB4uqlOAnz53/W56+F5mtExcpS7h5Z
5UE6E2mxCtJHjpZaNtVa2/jychEl8nSKG76SXzttAXyySwdMa0+VF1wZZdb0XcjJ
Ulsex2+R6zahJoAZOpG1eoLZZ7c1WuVHscfQtgBDSZFmeadb7+mIIYEqFOSgKr0N
C11evtqhnVLM15RYp+RQz9lgRu/lNDiUmMGHp8Odv6H3v52Mj/2+VVzA0VXw45y+
Br3kxHKBIPue6B1LJcVa6eYPN3sCTCo10stvoni6mv2cnfIj30VqYTclxv+B3IrX
LzbL7GboJH5ZoB2a0KJE6/+bv54WS8lK2TLAVDr6HLPHka2gQUAh84Fvhb6G0BO6
n4mwHGRBX/41g+JZAG3SWN/Fxp0QSwX35Br7poE0PlU3Trrwx1eKFfTOsaJU7nCz
irI/2SdJgm9Y/S+ryQT6P++5K+d2uVYVKEqU0OkwlSWVl9iyTb19D4Ru4SteAYtB
FcEsiRpQi0+L6/YmgPo3ZYy7hLLWfKYis1WxugURGV4Xoq+vg8Pj8nz88/ZrmJ/b
Z/VzbY+aJ1rVqWyCvWPzVMx+EsS4JCrVp4yoW115cOzcFnQKvMc5t2yURREsci4j
EV3u4uPoi1pOmkoxXJy9D2p4YukxVACuyyiWmVj7CcIgR769GaThhGO2cKu5+cuk
LXA2/LqjGaRw9wvyp4PgLL5kMrO0k5me5RY2WGp3ptrZucbL3ws/LH6Z+ycvE2x+
ktpJznFfJrnC9kZixFa3A7yGIJXf6POzb07TttWoCjLXA6svsJRINYVVpp7BGrQv
NvA/cZGhcp4L2kkLVC7Nj868oS/rpIgrQ1EfqbF+/W2ytLsfaIT7gSGJMyFhuQA6
nbOilpTjzdKT3dtuPe5f6BHaFCRdCV9d4tkGfKeBXxQhsUMnCyFvo3S/RQPZiWVD
Z94lyumGc+/E7xoG9IjXP8AE09TKpD46WiZr1bI+4L+Bd6KwTZehLBU8AHHGwSvL
CDYYNVdxCrcmC/opwJh69+ZRyuDs+3KVN/nkF+TYih4n+GROn3UULlXdcwrrXoR8
hzlEdhcY+zzwDdw62e/K9/qTwa8ZN+GGkSgtOxhkjyXIEqZiX4zmTju+jTXBQDSV
7oTI2l2P507YBSxk4gNPGKTS9Zwr26HcHVHB9aTgL69cEceWqjz5LXMA1wTqlv6F
Mq3AlT62z5T9FdZh9YDKNIuI3TONmaa5bbASAMjcysX9rtMPbQf/0MU6v/cmM4FE
1AkdOpxY7H1Ls3fLAcmoVk0ie9BjVS0U4C+zQJh64HanX18PqB19McqX6Uw882fG
m9JZNgpm2PtAghh4LlQD1RJlL7bgpn1iqg/fxjrnzMv6yTQaWJCAfvaYDtxh0KQ+
wtM+n2Y858PiHqBNxKZTK9zIy7QhdXtYMpA62PZyQrIbCcGlioFpu1Il26wqrdK6
IOP+rl///bkZc1G7rjOkQLbzCgmi3RIg5aPc6FX9OF4k8iOP+xB1tQco1i2cJQpJ
AqExHHpM05NHXEfylTLMsg4DJTtxHTSwK0DlI/YZ8Arczu9g90v53oHDlEYxlbxW
Od9QMi7XnfkzMdnA7PZkdAXJRtjbnQfTAhNKpRa1s/dkKHpCBusBhkmj8MKO3zn9
TGabISCPGYE/lm4iSuKUfpt/QY9rhCM+1FL+VgxlcO2Cdq7ghxWUIXDtjk32RUL4
t6C1tqcQzA1utl+42te16giGoZHU5E9kFObfRzSCnjZWMwQR+0JvldXCXgg0rkHO
dc1egEnoZTwwNbYdjTdVEvLz4o7sP01AkulPLDzyRYq6jDelkiYSl98UQV9PoAX6
CzMF3Ibfz+fifFzoyZbAIxbTLIhBb8d/vtzaBBhPjotGWSBrc6v5As1DKOGsYEei
a+Yf+DYAMC+OD56yhj8F1PK/mCfOkXbmkiYRqI8R2LZZLvS6pQYGMnOOWlUK2+tj
ba+L/rySr4dbNZKVyC+2p/CZ12zZ28PmmijUM+wWVQk8zGomLtd05ZV5WVgdI8I4
veK0S8+W3XizNOZXILJSYEOrzSaKE+jdhbdAsJSZs84ZV4wZKVptETCaSqbB3aqs
6JlKOqtKWzKgtrQAftcXu5jyxTcsqZqgCw0LxRT1dm5+U2SishfUPqDoUrRNdpS1
7yo7y4Njg7aZidZjSEDqaQE6qnMn2GiUvmFmRyFSwcStNoS+5gT9vsj0oB53ZmYX
wS5yTrF7A566CVP9hS1/0oLtLDy+bcaJMGYWOBg8q8xboOUlAQuA8np1MQQRWQh9
w8IZvp1Vo38e96c0uCnkYfseXGoCKVe6KNUl9S8iNE9puXxO2jJseXrBsYUrZ8BG
OS4cr4D3ZJeAsAc3cgWDmlehb3zbf5u0XuR55QccXYZsoYrz+l4dQBo+xsVDfW9+
VgMmAh/0RqDDf17fxuHCcbv40LbFjEuUqd2WXwzOm6aQcwCThJ/1EsZIG3IPdkbH
NTmLQFNCm7Xzh6hMgU7IB7v0o+22UD6I+0oPmd/nMjVJ/67WL1zM088A3RNi08og
K6MhF8XDZ5BNqPxhmbfwUwvQY7CHbfagpHqUR8VeT+7L1yMfXV6tiVPeLkc830sZ
/ZgSSswuBJJwUcWCSkcRl+FoTZskxkdF40QyFTqcPm49PUyA3/2wf3V32A3Jcae6
tZVoJfvndqNvJkgWe4g+6RPTmnsskmuR1ZUTizpm+5we9w5vm5BkrXV7eAkoY4K0
GpUtr+AHgEwTDdlAmFlAVyUaXhJPtyDBWgUXF8RtQaObllc5yP05pCrrIE4bjyxM
3qgKeFbKhCh/XCQcHdUDnQWVaHzJjyaiZy2nGQJxRtVWK9JLJxcizn9lnHT+pBov
B+eIDWGBN79DEBAHMt1d9ZyQors3awgTiVaELj3ALdCYF6bJbmEYO8y8TvqGwHP4
6h3hpDGBjm0rlD3MoNWf9pF9hbjrqAv73/fe/XH9L2ue2Oq5kXhA/FCEGUPYQinU
J3GX7vXyES37xDEQSEr66X2ScBNpJ0VrlwQTgTkkzFh/rOTC4MEERBgguWIRl2Q0
2i/jpFbMorhxvxmZmpYwL0zGlK1/DeEl93L1uDMzR2yueVKWBbl+5a9cW1gGVUxa
kDuTKupFHFg2hCNKxLp/pSROi+lJdudf6/jXjjn8PN5jtFoYDTJQBNPiwbdPrMyg
LCu+nhbZ0K5jBHBkhjWgN/NXNEhugyN4P6uayJNvx+mDeMMQ6TRd/0qk36lXl0mz
m4NuzljAq/povifMO78EiiLFXU7MrrtEgM2Ax5PwfuAojCnW4kwYrZLQ2hEH9B+j
9P2zUo2eKJxg3MosQ00OmePCjbSvIYda8r7ujewbu36Y4kSCUEExlgVKu2sLALjh
gHCtNpDHW6JBN1O5012oxrnjgw7rzs28HUUu6mDh8qJMSnaCDuk8I7wZMhdkVAjz
NmO6NZCriEWz9HJR+H7+iiueEtQiQFIWaON8PMMKgshsDJGANsKfdnWEDVqmk194
Q+52eL2jumvmBf46PPZdYa78PixMwfpMCuWTfzbKcvUui/ucc0Mmbo4Y1Jo3tWxm
4njjqwyZWWykgzqmPqWlG+sXrtqz/VpWT9WHyJR6xeO0NjF9XUa0SzcLB1xkq5Re
KPxJ0pvi1PGcY5fwf7rX3QGgdDPDhHODJYNTkw1djgpr5fkA0SzHbeIcLNBAJVod
RM2HM7zobL25wChwKPTDjcjH72cwAkUdGUhoL2gV3bx/UZ+8dGLfTBkfZHPzubQ5
DS7TQT7nKM81RGUFuFvb7LrBHOb6U4cuVX5sG6jjqQ8RtrVmtwRfgoBQ9iZNP1Zu
AplMO1pCkIZ/yXKrnxGC2XK3wTRbq8WusgpsjuF5IkBQMGthf0c4e+vNBPayg9Y1
K+YTwshy6WAU2NttzkLxRRRiUBhUma1Zj0F/oGNLCXf1zr0N6C2qnkw4p+O+BBhz
sO2eFLTJpKgCjz7A/buP4WnKFbuF1JzRbY+y0X0llbhw3hD8MoMafNjtv9Euj4dk
K1jwZV86VLD1O4ZaIUvvS3Dx0PuKrBIOq2Vs12QR/6D7X0kSNl+3AjYWfzBOBjaP
+PL5DtdG2Xsca+F96oT8J5nN3juvdBlpU6a1mSPVNqKMRJVPCvhru7iO0auL1tPM
Y1nUMWKwoC/ABH+YxRNCXtOcvJFraC2hX623Gb8lF9dWWqNQ3q768GBBySAwMKSJ
YJSWExXc6g5da2V0uAXND9SXLzmw2J4pi0JQaQ5ELtEIXov0y/lk9mJtg5E7Zhk1
UdjesZnDnS1ZgKjJn+yqnIoEEnMHUOMMATiUEW5uz8RIMi9lfqmmeihz8zXwF/C6
Hy3dvBVOJ9EU7St2py5iujEabHJC7GJlbcYzF3plRCH8EqP/AdmiKY0CuFqwRxtQ
/0lf0m270RULbj3/awQAivkiGfrU2P+BRM2zxZDRgVgDAZN8yA7Ln/gDvztw0SSG
Q/lKsJxOk4q+6YAMfmSiSoIJfwFIdsGYEeOYJJGIdtqHcAipXgGpZufq1fpzD+AT
BJyLUZFUyTDPH5eoVyJoEQ0EwZl8vf9Fzr3JrcHKzs8p2Fj78apOsnnjK5lVqqbu
3SMHeqYlyeLssnCU1pu/zOvcnFW4eCepnzOj3hCbXJka51Q+h3/Wm79AN2gAukJ9
LT7ZRi/9t1ibotYFE/W9vixhHY1yNBw/oWpA5ezEJYHLJRPNexX5/6c85cLR38wE
GnI3FKqDu5X4nLnD8OihCkRSOHnPOQbsOLiovjIn/BpkhBgtMk2O66hl6BumHq2q
r0qPDrLTTreboVSYXZxMuXBbDN+QmKk88p+QVXlsYjOVd3A7ZkhoS48yHXMz/S9/
7dknr0Bhn5/LdJ4NYA6vHpMtPizEZNlYHQgQmJzkPJl8eGZnAyBRRV2xnigjLoLX
Dw66sNJ91TB4n8p64CoJEnNQ/ZWgMuT73EwwOOtzP9zyX5MfHBeGoiADmwF1gp/D
33htFb5yUIZA7ITUH0JD3syRLn1KNcIkqZ3QV90WtpVN7YvR6+vl+ZQpO2Wh4x0S
SxEOBWDLMaG0jYnKUo3PU2gOQ0Pi8CTn5O0V0xfP1pxyO1DFvKQS8kV5oH2r4GRE
BXIW8odbbVM+eq3vKbNst6hIxyqf/zrsXi/hkjsfxmBgSLuZ769fSTvdxPIHvqoJ
ml9TeJVJNQBdpW9R8XK/69Ra2qAxoc6COAqh3/deY1w5fxUoMEW3bL8Q0sjELSot
fbpotVFl2cd7rfVek5L8kSxwSr92gmhaHw+YYeZLgJH92xLvulTYFcCN8NQkoUrl
XnRwz4FvPq5jGEgpqCxfJYabEjZqzQ1htjSDoARaK+WI6Cep6fGr8U2VqkkFo5Py
01zA0wdGpsW56NwEvJ5sXuPVXZW9ToWDG8gPaRGrk69ACCK3PBfwA0Dg5BJ+zi2+
mrKazDNQoMrE2a2qH/9vkA==
`pragma protect end_protected
    /* 
    * Instantiate the cfg for master only 
    * Enable timer only for master bus tracer
    */
    pa_cfg_xactor  #(
        .ENABLE_TIMER    (IS_MASTER)
    ) cfg (
        .i_clk              (i_clk),
        .i_rstn             (i_rstn),
        .o_enable           (r_pkt_enable),
        .o_connect          (/* open */)
    );
    
endmodule  
  
`pragma protect begin_protected
`pragma protect author = "MED"
`pragma protect author_info = "VirtuaLAB"
`pragma protect encrypt_agent = "RTLC VELOCE", encrypt_agent_info = "1.5"
`pragma protect key_keyowner = "Mentor Graphics Corporation"
`pragma protect key_keyname =  "MGC-VERIF-SIM-RSA-1"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype =  "base64")
`pragma protect key_block
JPKZQTCF3TfLqKFKk4Wd8RlI/rtSBtUtGuP1MrDj7XQEl1wRK41iOv4AuAOr+eE+
KbE0QozHU34qAwEiIl94n7a05PCBLJNHLG0HxCU6MBXHFwQgIqafwvIezaou4HjU
cq3jzfK+5Wd0MXcL7MVyXziXIAHCR/3cAMV8LXHCYT4=
`pragma protect key_keyowner = "Mentor Graphics Corporation"
`pragma protect key_keyname =  "MGC-VELOCE-RSA"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype =  "base64")
`pragma protect key_block
q3q29jdPOgbCD7Pl0tBf4EjaZEndinlwexCr88vKEE7lCBPrQZ13y8FQKofAUvcv
tY1/Suhb1fVK6T9Trpg92/4V4LqVFMrwjBL0Mpw3icsexgzsyiisJrAZuzQWLd9F
lOujaETbS5rNWxLmfFift2/ml/rVSzQB004dMVcYjZs=
`pragma protect data_method =  "aes128-cbc"
`pragma protect encoding = ( enctype =  "base64" )
`pragma protect data_block
XMfHdmFmTqCWCArz8t/U6yfAiJScEAjuGqu4PUJ63IiAjVfMXfG80FZYvube4Epu
niwcLmCXTHJpSJZ6lKzfvDnN5C90g/llvTA7PfM7Wulij5+xCmfFTiV9vD+R5OKx
E/Whmjb88bMgJWjQrFEnZ8fTnXOA/bD0DQl34Iku5uokmA7N+r5ui123tEhPtdYG
KtUUWyV91ryRGLbm4L9EyqHhY12H4zs9mCjbXtXweACDdyc+yyhVU/voEYVssCJt
Xq9fqSYkDkTqWSlTxmxGk3geXMhr9+i8vJxB9YSNEAoWJPth0nwIbVn/1Pn2tvsJ
Aexg7K+isOoqJqHoeUlnkQmiG1V/+y6CokfGISrVmXCEl0TYZjJzF0UjDcJKFtHF
NG84b6jlKZQuBQ4tR5X8SwshUGjIZ0/+ZgqPg3vjVDEyN9YnahI62KBirRTqVXc8
l7JOplLM8zgJc6n80OI8v3VsF4B70sXaVWLE5N5OhCys4rzgXnTFivIY+zff5/A8
R5Dul/gaIzvaSowmFox5mGTY3NInM8SqP+CX4W3gpRIt2BrJu53sD1apzPzdXVuz
cZQpnhpX1Y4c/+D+bVR38IaFyFpLjOQrtPWfFDdHgVc40i25iiLQBFkEJL9yyZk/
G9XORAnj7xbwtu4P8U30LnJg9izbOjsMCR2kaK4OIbGRpISStRjxrjTc/WC0E4Eg
IsWoVByjzchiZhOhhhEyANcAQ3JMxdssRTPXyftCaoYJn4rJ/D9DVSv7ZYaMwqv4
IUlonKHdYf6d/Z+eC75CxvYK1MppEGSAlODU4bWeMVXMsZBs/COOZYT9AqMorZ5b
Lxas8OuskxjuLUEEDAj/9/NXL4eNn28mZFJSsrimLr549x4oByGr8gu+D2SDt4ut
AryYPkiULmBFLQPXTPiof3sn0hbE/SygsbfCUbg732wHWrZ2l9z4D1tkdqLZMdV2
6VFhyRk6exuoZi+Q6EHsy0vjAkAK9RDmfe6BPp1GGxnQDQ1o6QZkDIIVgKxuD5ea
dAJ+Pqp3U6G4LUwXzC5ZiMdVZ41GHcTriZojBW+qaq4fiLjZQTHvnfVKhBb7sYa/
8cwkoyLWnx0RfOPL2dknOrWBQJtoKZaQfjzBlYbXn+wOEb5BY7ZDyrFq2hjMuWnD
CR5H8IkQMnMe13EVlC2zFB5dTZbOxpVSASwIoxg76+fH5l9YKbp6b1nbT+YZwv3N
CA91i8FoV2+19ZSmQbcYRqrmnvW6cEmQZSBycOnu0CXU+vl6l/xK4fc8VaNJSWi7
RS5eYjo46GZsvMX8ga7N8gnLGVyOt67d2igjzZFKAteOVBa7Mbc9nJ+9w1yTT8+u
jPm38I8ol0DbQJf9QjrY/pKHmvbUw1glcUcWI6rURTd0YFCuWRBHSr+NOaQ/oS1t
dqhk0B50oOLb+vZ3dgo8jzinNKfrg4GOgktahFgsEf9rBEciktLKFRmG4EPIeC4C
9wWngc77ABerlUSjJ9KHPHdWjdl3mQYSRBVYVMsFD4ZmQMkL2jYMhFDlrkrl+6pk
Hg1Cf6cqH7s31ABfJ4wvuLCVnDg/RuQ7RT2k23f4EsRyxSUVhSnhhlsy3BLqMSqK
rW2PYbND+KoelQhl/OFTF+eimJY1K9/IAxd3WO5QZOprKtFDZEE+xsLG6bBqMYBJ
cmQiUDIY9T/zlM++q/GdrNlYtn+olJtbZlsiArOZkJMX4DRWDrdwudGTR4tZGAe9
dTO5sV220SMqIxC5Fr8+D2FeLh8k03GOa7/UbZlZpiKqkTHW8iuKXc9xXMxootCG
4RThjxdVLbkiFOpNaKTh2lgnLyEZITn4bIxHkHTv5moh/FdRR7FciX+3HY8OfeL4
/ia8S3m8KZO0It+uOqDpfRvd5pZJvkX3t+75+NQ4nWmGLwO2C+IH+2xGWOPs+fFn
qoik/GL0P4WRCZLMIKDTM59MylaGBV3sykYwCnfpMbxsKQYgHmYpjI1sE9sJN3pB
xjoLHa2HKIVKBZmvh2bGn5Cku8x4J4APujeG8dmlcMWOVoU23ZheN9/qK8EKDNzv
H5wGQ7W4zSVbi+6ei0ATdq0VOKdl5/jv0BDEKUePm03YnucRp4BOR048iw6XDk8A
zQGW2GI6R0VWfAEtFv7k89O/LhAkDecr4rQ+1d7RhE4QQqocse+qnhQ3yEu6/9HM
yYgPnTs5ePzJih7V3rZozHvC5HQpUU+YlGJlJel3AHsq9mWZKOqlqSBhGZJQQWFu
2NpopzF5X+042MGUk9Q4RA==
`pragma protect end_protected
    /******************************************************************************
    * DPI Imports/Exports
    ******************************************************************************/
    import "DPI-C" context function void on_pa_cfg_timer_fire();
    import "DPI-C" context function void on_pa_capture_changed(input bit [EXPORT_DPI_BITS-1:0] old_enable_vector,
                                                               input bit [EXPORT_DPI_BITS-1:0] new_enable_vector);
    import "DPI-C" context function void on_pa_finish(output bit [31:0] dummy);
    export "DPI-C" function pa_cfg_trigger;
`pragma protect begin_protected
`pragma protect author = "MED"
`pragma protect author_info = "VirtuaLAB"
`pragma protect encrypt_agent = "RTLC VELOCE", encrypt_agent_info = "1.5"
`pragma protect key_keyowner = "Mentor Graphics Corporation"
`pragma protect key_keyname =  "MGC-VERIF-SIM-RSA-1"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype =  "base64")
`pragma protect key_block
QtW1MRkLwNTqo5MJ41fAobVNG5jiUyzAzaZEARgoB5JgMmoCOLcG4sGb1Ix2x6kX
/1lw2v9B94aUU1D0DhlXC62NpWBUcU83Zh4t9p/CtCy7IqPK1eGdhyxUZtY6wrAM
Jov5n5foeRlrxIhtg3QQZaaivqACTOZyoa06sDzm4xg=
`pragma protect key_keyowner = "Mentor Graphics Corporation"
`pragma protect key_keyname =  "MGC-VELOCE-RSA"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype =  "base64")
`pragma protect key_block
fQ+0B9atuCCMbOr8KHjPg9nt+P/pv12GWvDczxjkBlnQeN3i2ZNEhL1uCEeolP/s
Veqp0jXuXuMBl2enaR5x4QEZ0ax/s6SY5JzBSbuPM4WhfoeXLZ79UqMS9rrF+cRU
n4+B7/1ohyot76xZktrtpLUW/jIgAM7utuCNjbW1fSQ=
`pragma protect data_method =  "aes128-cbc"
`pragma protect encoding = ( enctype =  "base64" )
`pragma protect data_block
JMi6Wy7uVW315RtwN0zkuMWfEqnIRikfIDzeYp1docLA1K4VabbcmLW22QGKPzRu
wHYQLKb6mPtyQ6avHAi84+zgbIQldgC+mSXy5fpHbbGLkjH6MILDOOoVBkKRjsA3
koqNyyvF+GH8qh1DuJT5xXAvm1IQTblhtTZ/PrNECkcZZpZrnA09krt9uwbduxYX
DtAPYLlxUqchktzQnYQBTETbhVYfs19OrAXmo1FRbVuYAdfGpBkCvMsBzWIqSXD5
ZlU9BKf8ic7Gu2Cyb+7eOt20Z64MGKr2yRSOjOjMEqVmAK9t2z7OucoK5Bjw9PTb
/7W5s5YMtXU0w6D2dbtL2dLwyugXMjJ20Cco8QpaPuMeJ87rMK4g9hKiWcwPvgRT
ckHtMbK057AOfif1zvTTrXdJl5bh85xXdTjcREZG5p8RDTSybrgirtd/1Prc8BEY
UNWb69/Odi3dX5kC4VuwQ2eAiuyUAyTD0ivNSPX+FfuC1UNb13/yvRdzGZ+lO+wR
NAFJc239PDKqU5uuiLXXPIwkrby29X4Y470+9K/eFc6zAHtkfibQkTC+Z7CptHcZ
PCyN1PPEKgjA6MqakbFShBEMxYnGqEAfiDvdxvIVkt/GMakE/XbSyviGqe1bVSdl
fGL+DVvKqHc0JMFIxKDEq55iPFpZdI+ylr00XuABH/cd3PG6U9b4wuoKlDva6hWp
zaLCm8KzpLN3RP/34egKmUy9SfrxIGgSJnDDDdxf0iOzDD+e/dJv68goEd0i2NMx
HR7ZUUImwzDWAwlBDQYQksarmsCDGpMHT0rsaqwwuR0eQE9jsPqBPoZQ5BFu2vm/
QDAYN50Evh0Bc0i4SxTY5+UoYO3r4n0LI+PtWU3tpCu+I4bllovPy8oA56Ntnsnn
qxrp2ybT/EufTSdtCCNv3LGWhVRERk/kDtp5ZnGN2X0q6JFqYDNFE7Qul0nklPKo
BiP7UTTokzWoq9LpdQ18eNUi5ur8bWobbPZEasHUkxmY4GcXI2Ut5GmCeMfDEQ4r
nZwG6Zv5HRllagEbYc5Nwe7U5imcNZaYG8cwTp4I/RnsLJ3CglFnj4boApNDKa0p
MlAuMZYTOYfbzHKj1WZHmkAZsNbiUlkR/95LMw660O1yCou8DKHudEBMz4TgMM/C
LdHu1DKpRRukw9pV1vsXap3qfpZiam3U4u+aCEBKrrbzaQJ6e1uzaSRrkouPO82b
sSSmqNrQfc1AEHYUTG8pzKzm3IqeFbrXaEfJLUXjH6sAOEuwY1b1k5SJUxShnu7J
qpy1BJStUbK6Fwnd0qb2Qe95GNW20ucOp8Ed5SgmZh5KBBj36lDZUVkZbuQAS/2P
w+vGnIVmYcioW2d71IJi1TrhCGAgsAja/g1tjdqA7ZJfPzIl5JFqUOZlvhyvazg4
MPv5D5yoHo+TogJHu9MlsrmyrUsMcB7gkpzM4pVF70YpUef0KqKeGuTy2aUPPiOz
J0z8J4iJniPQAXnGM8gL+KUVOgcR1WUqUqx3AaiOGvrOXVKjhq7qWWbEZMQIIiH7
l3V7vQ8c52/RPT7kJcTdUpASJXhpSWnvzsUq9QHSzoB1Lx6Tq4kws4WGYt1voU4f
UpbJlu0D16xR8CUwAyXxRsD7zheE0Ny1BTYztV1JDycdf4Eg9D5dN525JJnvDMS0
nX4BzrkSKEc0JPibmBr9V7Klhjj45YQJ2iXi6nDhYW0QneRsIfx41UV98n1EqlZi
oLxobkYE4WLFMDSJlKbKrcloFumYU9pbqjNatzz+HG6kcPTGiARtGM2X74z2d6TX
myJEhwY3c3pIAJbgIoCyDKgg/nPQTYXSNVmaaomQAkpAJC9ywX/tcwODf6OKda7M
vrs8JIsiLhT9tMRkb0DS931VdC8ni2przRDsTcJ6K1k6LIt7mfEbA4dyJGmjCZh+
28X7KGpcYvwxqfg1gESKaJR/vvbz4ArQYCan8g/r70uCxrNYRfuVoB6s11bM58DF
C/iZ55MtwEjZeByqIvTP/sgZ1atafHEv1QZ0nh0Rb3/MzSqiwUtfpy4Lf1iJWvr4
NA9If1r0Z5gbpg/l48PrnJbCGqeOoIRzqvhpu9fiz1d3+yLylxj0H9nKkPkNTxkc
zjgaCSII1G9KzlqmgeCWGXMGLkpNqfq8pm2+cD7cwQgJPTKfcW6MKi4rzHUVIyM/
b5mVpUXzise6Gk3oKzq5d8vs0lDHQhnFvcD4laVSpAKdrEYw6JSoFU+38TafRxZ2
yDR3aqwAVa2EeIzxRpl0ZYjABktqvZ16wpOexDc36baACe56BN0DWtf5ahFSmRz1
zjlProaQsBNV4/x/TVcAF8+HPqyqPPHo4+96F19/SVuG8LZMgy3dkJ0As2pFCOcy
FzWFZkYW005yJHWekSN/8RoggLe3aNB4ZfHTd0VYdnVy0kPj8mJWNvkETNXqVsml
RWeFKiwJ68Eu5d/DDLoweP3zxFEzBY4Z0kpHnTR6PmxBlUjEs9OE8jn7/n5/2k5T
7ZdyD3kE2xvitPkbaEVXKmQ9rVYKbA/8sdAtv8aSqtrkN9j3GfSTxGrLAdeofoHP
6hBra6LEUzkAMbyC16ByIurtCBKctGLei2ZSvve/UjP/mZ1JfPezK9nsVQvXRAnv
WSeU4WUUA+nJwLK9AC90X/ly9qLq3i9HJlEPFGl7dOlNuXEW+cLg4Dj3D94SXEBp
jAkxAKMAxkDwfwaGjgvuUaBfY/cdV14HzEOLod1W+nNwgeXtgAjC6R1Olb0Rx5Wi
9AwYlHIgP8Mlz/l19RbbaBSKs1JLOZbctx+Jg6+JsLOTFpAbCetccMWyC811SvUD
Rv9sJZe/GVmoZr20bR34HSXCTyiN4GxYWWY3H6qKFyING5p0h5LlDZX6+lBf8DA+
3Ctw3HNAWTMiidB2sEBM25sjOo28rX0dY/WhmBh6oaekiWhSrhVF+UnwJVJ6WBnI
Ui64+jpzPQO3+SPOX8T6xGNz6WBQAF4TchqZWnb6soXa1JNlFd8R/bDW7CLY6zm2
uO4Bt7p+3xrD22niU/9A/JVqTqXSb5wwtmmyRiqMrN9ActX2mz+0WmjZuFNapr6y
asCRUAOgkzKv1B6UnvuNwl9wiHAcb8Jj3UsSCo9tL446N73HfnU22tpk8LnZfb+2
qRX3G4F4imqbIUhOlFNZpWzZzzPtpzWuop2LluDxkPTCtWlfI7/xVrAqofNT1451
s5yMa4/JWGkkLIBKAcbRoEllB85U5gQxuFhe9fcBJ3zf4MNbkL77nmH8h8ueMZHZ
bcH6QJIIlXzBTRorhs2RT7wdWJF6mWYYZjv1KX8jYoTq5oX1AV/yp//3XQE4iwXC
BLq5Jq1yvhyZu11pIaOvIFxSyn8Ffn9SWsEORB+DC6tnxBJdWVm9ZPQAtNe+RfbA
JSR9P0ZC/zWd+2d30Jtbngp47DY/BkC8uaaGPrjHJ1NUH7JzyDNqnqPcEP8/n/GT
MZ3XgjKwEuhhbyneFpXiVUR9H0NaVRsnRa9+P6sP1UEKl/kS2Y5707yPo6VEj7yW
ELDGYtT4UpbNcK1uPInIwRsShuGj0OVst26gqAynpSJTkThoewZVzWgZ/XHQf5Od
g99ePBztRGirhoq8uAPStR2wd82oxLc+AMx7veZj2nG4C4nVdsgKPg1TnLOvPkjo
AsDUDW8HMt2xfShe4xx5lecECxjHDFaLS9+bIHDNCPI0LLkBKCljkosod6JM8Wfy
GdkH3Ys+7AihYUxF3LhYGEpbHNR7GzyCHnU7p1SCIApyk+FWgyfuiFDWZdknj4JW
ucFrcNZXuELGXSSf5s9TZYbCVZs6W4VOcvbG5H9w+DMRc58dS+vA8R6HSonByzrq
atzeTKg9vh94wlsm7l+hMBsCCXl3fCQCFkfCi0UWKt2nmW3tjQWAfHnkIp6B+c9w
62BY9Zlg6daoVnV6kR5nl70FZATCSuTCbKMaUs/uV6qmPtroWAbRb3SIQPzAfnjV
EsD7DD0ar6iEuFzZfwSX52H//w/+W0nbFdn78egQydN5mw0K8wc5qV43vHRn/m7T
lnLdYpFybKWmey3mBD1UzJpp+cd1Pu4KTuZECsX47I6kz1Ot9e6Bh2jTSlSrS5AS
j3jqelarVO2sdRJIheZU6/Qd4xaFnjNUipjvz+3lapMHCkTY14XBH7xLU/vmX0W/
Tyt+s0nbjNFmS/A4vH5G3SLTpyDs+ma294tWd6M5RwxraoeBHauKynCEsCZfYpzH
/7F6aP6GErVvXLhhF4W3itDYDLMZWkf1LLKzszVcgQKF8Dr8bAPq+G/Ir2gXsBHT
yGToHSh8EkUid9sWrJLSBr5Uz7KJ7dD5bN7RhCbvYl8o05x/ePAXcqmbQeV+8Qzt
vlgfDS4FSV30ZoaRALcMvYrLveodKKqjmPeOr4tbn2t/yjHT0nD0b/eCwOzgEsfP
XT+lKBDwosZuNCE0FV8Y1R4H2kM0Ar2bVvKDdFSvSBWrxoAz40jBR2sBuX8ZcXbX
2O7JflGmYLMYYfGu3Aw+G58A0qiDqVRjVKdol7+Uw/S5JUr41bQQNUrmd26dvso/
WxHJk0TjaFNqiHOT6M6cbXwtiIFJwycPM6voQLaZo5rq1pvuzU1qi3TWJlfKkJrI
29bQI43EPQxOO7VvNZvOr7rUfg+PCiM5tgvZNm9DmSYyU2GANlLdZKp49iOLCVGQ
2EBOdffkXnvxR+Ez23EM6jCvfAgVp9Z4fGgoX0bsL82oVlI9Is/qLaZOGv0+ORhC
x19S/tGWiZ4214vJlvs6JyADjSvVmLVcxeiu2hbeG+UL1pdS/lWfADkCOsuRqv3f
BXOZB7N59548Z35Q2BcFHLoMp+HqoE9LJUlQI3FspejVF5K0v314mVt3DjeEmeCU
SUW8KDkeaq0SkPT1SAjnD/Irv7NsnGD1ivYVY3jPP4UDd3yqqjXUWOXX1O2tO/Gk
4LlsRKLJxQwijZwHmEA/tDsh1eTP4Xi5wuhd0az5HwKtlhG6E8eXFhg/icek3cM8
f07GBNL6YCsUgYo1TFoB8l4BhCCEvqXz7lraT9Z4hk/jIDt8UFmB8IWLV9hWfbMn
uJnurnzYPHH5V8jb/6+zTRyfQRZOkViOHS2P4u0yTi6oNjgkP4Nyf4hOWLcRjJAd
BRS1QPWrMmBB60htBVUbTdZEHOUFf4bFI73F3zULURtD0hTp70PVUL0BCCWyRdSw
RZmaiVkcBdoFwd2jpVixh2vtpNIvNDMtz7ZVuFzQ73h5GiA7SxnoTFvcanE/615E
/rzxjJRucgaVnYsldMpyYB2vOb3a1bSVNPOg9prD+gu1ycRIXujBsOkMZYKl3c0f
eSZ/kxHfs9XennFZjVOB2Dhhd9cEvRH+0jA1diGLk22kaFs/OIlCu0wA0vJIhiUV
p+mlprWD0r4GenhY+CdCvHcjjW2t9vu8Sl1i0sxSsGYTiVDaThIzTMtFi2FouFYO
iQwS7TQIxUPPjuN+yi1B4A==
`pragma protect end_protected
  
